-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b80c4",
             1 => x"800b0b0b",
             2 => x"80ca9504",
             3 => x"ffffffff",
             4 => x"ffffffff",
             5 => x"ffffffff",
             6 => x"ffffffff",
             7 => x"ffffffff",
             8 => x"0b0b80c4",
             9 => x"80040b0b",
            10 => x"80c48504",
            11 => x"0b0b80c4",
            12 => x"95040b0b",
            13 => x"80c4a504",
            14 => x"0b0b80c4",
            15 => x"b5040b0b",
            16 => x"80c4c504",
            17 => x"0b0b80c4",
            18 => x"d5040b0b",
            19 => x"80c4e504",
            20 => x"0b0b80c4",
            21 => x"f5040b0b",
            22 => x"80c58504",
            23 => x"0b0b80c5",
            24 => x"95040b0b",
            25 => x"80c5a504",
            26 => x"0b0b80c5",
            27 => x"b5040b0b",
            28 => x"80c5c504",
            29 => x"0b0b80c5",
            30 => x"d5040b0b",
            31 => x"80c5e504",
            32 => x"0b0b80c5",
            33 => x"f5040b0b",
            34 => x"80c68504",
            35 => x"0b0b80c6",
            36 => x"95040b0b",
            37 => x"80c6a504",
            38 => x"0b0b80c6",
            39 => x"b5040b0b",
            40 => x"80c6c504",
            41 => x"0b0b80c6",
            42 => x"d5040b0b",
            43 => x"80c6e504",
            44 => x"0b0b80c6",
            45 => x"f5040b0b",
            46 => x"80c78504",
            47 => x"0b0b80c7",
            48 => x"95040b0b",
            49 => x"80c7a504",
            50 => x"0b0b80c7",
            51 => x"b5040b0b",
            52 => x"80c7c504",
            53 => x"0b0b80c7",
            54 => x"d5040b0b",
            55 => x"80c7e504",
            56 => x"0b0b80c7",
            57 => x"f5040b0b",
            58 => x"80c88504",
            59 => x"0b0b80c8",
            60 => x"95040b0b",
            61 => x"80c8a504",
            62 => x"0b0b80c8",
            63 => x"b5040b0b",
            64 => x"80c8c504",
            65 => x"0b0b80c8",
            66 => x"d5040b0b",
            67 => x"80c8e504",
            68 => x"0b0b80c8",
            69 => x"f5040b0b",
            70 => x"80c98504",
            71 => x"0b0b80c9",
            72 => x"95040b0b",
            73 => x"80c9a504",
            74 => x"0b0b80c9",
            75 => x"b5040b0b",
            76 => x"80c9c504",
            77 => x"0b0b80c9",
            78 => x"d5040b0b",
            79 => x"80c9e504",
            80 => x"0b0b80c9",
            81 => x"f5040b0b",
            82 => x"80ca8504",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"00000000",
            89 => x"00000000",
            90 => x"00000000",
            91 => x"00000000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"00000000",
            97 => x"00000000",
            98 => x"00000000",
            99 => x"00000000",
           100 => x"00000000",
           101 => x"00000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"00000000",
           105 => x"00000000",
           106 => x"00000000",
           107 => x"00000000",
           108 => x"00000000",
           109 => x"00000000",
           110 => x"00000000",
           111 => x"00000000",
           112 => x"00000000",
           113 => x"00000000",
           114 => x"00000000",
           115 => x"00000000",
           116 => x"00000000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"00000000",
           121 => x"00000000",
           122 => x"00000000",
           123 => x"00000000",
           124 => x"00000000",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"0080c480",
           129 => x"04828cf8",
           130 => x"0c80d4de",
           131 => x"2d828cf8",
           132 => x"08838090",
           133 => x"04828cf8",
           134 => x"0c80e1d3",
           135 => x"2d828cf8",
           136 => x"08838090",
           137 => x"04828cf8",
           138 => x"0c80e292",
           139 => x"2d828cf8",
           140 => x"08838090",
           141 => x"04828cf8",
           142 => x"0c80e2b0",
           143 => x"2d828cf8",
           144 => x"08838090",
           145 => x"04828cf8",
           146 => x"0c80e8ee",
           147 => x"2d828cf8",
           148 => x"08838090",
           149 => x"04828cf8",
           150 => x"0c80e9ec",
           151 => x"2d828cf8",
           152 => x"08838090",
           153 => x"04828cf8",
           154 => x"0c80e2d3",
           155 => x"2d828cf8",
           156 => x"08838090",
           157 => x"04828cf8",
           158 => x"0c80ea89",
           159 => x"2d828cf8",
           160 => x"08838090",
           161 => x"04828cf8",
           162 => x"0c80ebfb",
           163 => x"2d828cf8",
           164 => x"08838090",
           165 => x"04828cf8",
           166 => x"0c80e894",
           167 => x"2d828cf8",
           168 => x"08838090",
           169 => x"04828cf8",
           170 => x"0c80e8aa",
           171 => x"2d828cf8",
           172 => x"08838090",
           173 => x"04828cf8",
           174 => x"0c80e8ce",
           175 => x"2d828cf8",
           176 => x"08838090",
           177 => x"04828cf8",
           178 => x"0c80d6eb",
           179 => x"2d828cf8",
           180 => x"08838090",
           181 => x"04828cf8",
           182 => x"0c80d7bc",
           183 => x"2d828cf8",
           184 => x"08838090",
           185 => x"04828cf8",
           186 => x"0c80cfd8",
           187 => x"2d828cf8",
           188 => x"08838090",
           189 => x"04828cf8",
           190 => x"0c80d18d",
           191 => x"2d828cf8",
           192 => x"08838090",
           193 => x"04828cf8",
           194 => x"0c80d2c0",
           195 => x"2d828cf8",
           196 => x"08838090",
           197 => x"04828cf8",
           198 => x"0c819eb0",
           199 => x"2d828cf8",
           200 => x"08838090",
           201 => x"04828cf8",
           202 => x"0c81aba1",
           203 => x"2d828cf8",
           204 => x"08838090",
           205 => x"04828cf8",
           206 => x"0c81a395",
           207 => x"2d828cf8",
           208 => x"08838090",
           209 => x"04828cf8",
           210 => x"0c81a692",
           211 => x"2d828cf8",
           212 => x"08838090",
           213 => x"04828cf8",
           214 => x"0c81b0b0",
           215 => x"2d828cf8",
           216 => x"08838090",
           217 => x"04828cf8",
           218 => x"0c81b990",
           219 => x"2d828cf8",
           220 => x"08838090",
           221 => x"04828cf8",
           222 => x"0c81aa83",
           223 => x"2d828cf8",
           224 => x"08838090",
           225 => x"04828cf8",
           226 => x"0c81b3cf",
           227 => x"2d828cf8",
           228 => x"08838090",
           229 => x"04828cf8",
           230 => x"0c81b4ee",
           231 => x"2d828cf8",
           232 => x"08838090",
           233 => x"04828cf8",
           234 => x"0c81b58d",
           235 => x"2d828cf8",
           236 => x"08838090",
           237 => x"04828cf8",
           238 => x"0c81bcf7",
           239 => x"2d828cf8",
           240 => x"08838090",
           241 => x"04828cf8",
           242 => x"0c81badd",
           243 => x"2d828cf8",
           244 => x"08838090",
           245 => x"04828cf8",
           246 => x"0c81bfcb",
           247 => x"2d828cf8",
           248 => x"08838090",
           249 => x"04828cf8",
           250 => x"0c81b691",
           251 => x"2d828cf8",
           252 => x"08838090",
           253 => x"04828cf8",
           254 => x"0c81c2cb",
           255 => x"2d828cf8",
           256 => x"08838090",
           257 => x"04828cf8",
           258 => x"0c81c3cc",
           259 => x"2d828cf8",
           260 => x"08838090",
           261 => x"04828cf8",
           262 => x"0c81ac81",
           263 => x"2d828cf8",
           264 => x"08838090",
           265 => x"04828cf8",
           266 => x"0c81abda",
           267 => x"2d828cf8",
           268 => x"08838090",
           269 => x"04828cf8",
           270 => x"0c81ad85",
           271 => x"2d828cf8",
           272 => x"08838090",
           273 => x"04828cf8",
           274 => x"0c81b6e8",
           275 => x"2d828cf8",
           276 => x"08838090",
           277 => x"04828cf8",
           278 => x"0c81c4bd",
           279 => x"2d828cf8",
           280 => x"08838090",
           281 => x"04828cf8",
           282 => x"0c81c6c7",
           283 => x"2d828cf8",
           284 => x"08838090",
           285 => x"04828cf8",
           286 => x"0c81ca89",
           287 => x"2d828cf8",
           288 => x"08838090",
           289 => x"04828cf8",
           290 => x"0c819dcf",
           291 => x"2d828cf8",
           292 => x"08838090",
           293 => x"04828cf8",
           294 => x"0c81ccf5",
           295 => x"2d828cf8",
           296 => x"08838090",
           297 => x"04828cf8",
           298 => x"0c80ef8a",
           299 => x"2d828cf8",
           300 => x"08838090",
           301 => x"04828cf8",
           302 => x"0c80f0f4",
           303 => x"2d828cf8",
           304 => x"08838090",
           305 => x"04828cf8",
           306 => x"0c80f2d8",
           307 => x"2d828cf8",
           308 => x"08838090",
           309 => x"04828cf8",
           310 => x"0c80d081",
           311 => x"2d828cf8",
           312 => x"08838090",
           313 => x"04828cf8",
           314 => x"0c80d0e3",
           315 => x"2d828cf8",
           316 => x"08838090",
           317 => x"04828cf8",
           318 => x"0c80d3d0",
           319 => x"2d828cf8",
           320 => x"08838090",
           321 => x"04828cf8",
           322 => x"0c81daf2",
           323 => x"2d828cf8",
           324 => x"08838090",
           325 => x"04828cec",
           326 => x"7082a498",
           327 => x"278e3880",
           328 => x"71708405",
           329 => x"530c0b0b",
           330 => x"80ca9804",
           331 => x"80c48051",
           332 => x"81f3d704",
           333 => x"3c04828c",
           334 => x"f8080282",
           335 => x"8cf80cfd",
           336 => x"3d0d8053",
           337 => x"828cf808",
           338 => x"8c050852",
           339 => x"828cf808",
           340 => x"88050851",
           341 => x"80c53f82",
           342 => x"8cec0870",
           343 => x"828cec0c",
           344 => x"54853d0d",
           345 => x"828cf80c",
           346 => x"04828cf8",
           347 => x"0802828c",
           348 => x"f80cfd3d",
           349 => x"0d815382",
           350 => x"8cf8088c",
           351 => x"05085282",
           352 => x"8cf80888",
           353 => x"05085193",
           354 => x"3f828cec",
           355 => x"0870828c",
           356 => x"ec0c5485",
           357 => x"3d0d828c",
           358 => x"f80c0482",
           359 => x"8cf80802",
           360 => x"828cf80c",
           361 => x"fd3d0d81",
           362 => x"0b828cf8",
           363 => x"08fc050c",
           364 => x"800b828c",
           365 => x"f808f805",
           366 => x"0c828cf8",
           367 => x"088c0508",
           368 => x"828cf808",
           369 => x"88050827",
           370 => x"b938828c",
           371 => x"f808fc05",
           372 => x"08802eae",
           373 => x"38800b82",
           374 => x"8cf8088c",
           375 => x"050824a2",
           376 => x"38828cf8",
           377 => x"088c0508",
           378 => x"10828cf8",
           379 => x"088c050c",
           380 => x"828cf808",
           381 => x"fc050810",
           382 => x"828cf808",
           383 => x"fc050cff",
           384 => x"b839828c",
           385 => x"f808fc05",
           386 => x"08802e80",
           387 => x"e138828c",
           388 => x"f8088c05",
           389 => x"08828cf8",
           390 => x"08880508",
           391 => x"26ad3882",
           392 => x"8cf80888",
           393 => x"0508828c",
           394 => x"f8088c05",
           395 => x"0831828c",
           396 => x"f8088805",
           397 => x"0c828cf8",
           398 => x"08f80508",
           399 => x"828cf808",
           400 => x"fc050807",
           401 => x"828cf808",
           402 => x"f8050c82",
           403 => x"8cf808fc",
           404 => x"0508812a",
           405 => x"828cf808",
           406 => x"fc050c82",
           407 => x"8cf8088c",
           408 => x"0508812a",
           409 => x"828cf808",
           410 => x"8c050cff",
           411 => x"9539828c",
           412 => x"f8089005",
           413 => x"08802e93",
           414 => x"38828cf8",
           415 => x"08880508",
           416 => x"70828cf8",
           417 => x"08f4050c",
           418 => x"51913982",
           419 => x"8cf808f8",
           420 => x"05087082",
           421 => x"8cf808f4",
           422 => x"050c5182",
           423 => x"8cf808f4",
           424 => x"0508828c",
           425 => x"ec0c853d",
           426 => x"0d828cf8",
           427 => x"0c04fc3d",
           428 => x"0d767971",
           429 => x"028c059f",
           430 => x"05335755",
           431 => x"53558372",
           432 => x"278a3874",
           433 => x"83065170",
           434 => x"802ea438",
           435 => x"ff125271",
           436 => x"ff2e9338",
           437 => x"73737081",
           438 => x"055534ff",
           439 => x"125271ff",
           440 => x"2e098106",
           441 => x"ef387482",
           442 => x"8cec0c86",
           443 => x"3d0d0474",
           444 => x"74882b75",
           445 => x"07707190",
           446 => x"2b075154",
           447 => x"518f7227",
           448 => x"a5387271",
           449 => x"70840553",
           450 => x"0c727170",
           451 => x"8405530c",
           452 => x"72717084",
           453 => x"05530c72",
           454 => x"71708405",
           455 => x"530cf012",
           456 => x"52718f26",
           457 => x"dd388372",
           458 => x"27903872",
           459 => x"71708405",
           460 => x"530cfc12",
           461 => x"52718326",
           462 => x"f2387053",
           463 => x"ff8e39fb",
           464 => x"3d0d7779",
           465 => x"70720783",
           466 => x"06535452",
           467 => x"70933871",
           468 => x"73730854",
           469 => x"56547173",
           470 => x"082e80c6",
           471 => x"38737554",
           472 => x"52713370",
           473 => x"81ff0652",
           474 => x"5470802e",
           475 => x"9d387233",
           476 => x"5570752e",
           477 => x"09810695",
           478 => x"38811281",
           479 => x"14713370",
           480 => x"81ff0654",
           481 => x"56545270",
           482 => x"e5387233",
           483 => x"557381ff",
           484 => x"067581ff",
           485 => x"06717131",
           486 => x"828cec0c",
           487 => x"5252873d",
           488 => x"0d047109",
           489 => x"70f7fbfd",
           490 => x"ff140670",
           491 => x"f8848281",
           492 => x"80065151",
           493 => x"51709738",
           494 => x"84148416",
           495 => x"71085456",
           496 => x"54717508",
           497 => x"2edc3873",
           498 => x"755452ff",
           499 => x"9439800b",
           500 => x"828cec0c",
           501 => x"873d0d04",
           502 => x"fe3d0d80",
           503 => x"52835371",
           504 => x"882b5287",
           505 => x"863f828c",
           506 => x"ec0881ff",
           507 => x"067207ff",
           508 => x"14545272",
           509 => x"8025e838",
           510 => x"71828cec",
           511 => x"0c843d0d",
           512 => x"04fb3d0d",
           513 => x"77700870",
           514 => x"53535671",
           515 => x"802e80ca",
           516 => x"38713351",
           517 => x"70a02e09",
           518 => x"81068638",
           519 => x"811252f1",
           520 => x"39715384",
           521 => x"39811353",
           522 => x"80733370",
           523 => x"81ff0653",
           524 => x"555570a0",
           525 => x"2e833881",
           526 => x"5570802e",
           527 => x"843874e5",
           528 => x"387381ff",
           529 => x"065170a0",
           530 => x"2e098106",
           531 => x"88388073",
           532 => x"70810555",
           533 => x"3472760c",
           534 => x"71517082",
           535 => x"8cec0c87",
           536 => x"3d0d04fc",
           537 => x"3d0d7653",
           538 => x"7208802e",
           539 => x"9138863d",
           540 => x"fc055272",
           541 => x"519b843f",
           542 => x"828cec08",
           543 => x"85388053",
           544 => x"83397453",
           545 => x"72828cec",
           546 => x"0c863d0d",
           547 => x"04fc3d0d",
           548 => x"76821133",
           549 => x"ff055253",
           550 => x"8152708b",
           551 => x"26819838",
           552 => x"831333ff",
           553 => x"05518252",
           554 => x"709e2681",
           555 => x"8a388413",
           556 => x"33518352",
           557 => x"70972680",
           558 => x"fe388513",
           559 => x"33518452",
           560 => x"70bb2680",
           561 => x"f2388613",
           562 => x"33518552",
           563 => x"70bb2680",
           564 => x"e6388813",
           565 => x"22558652",
           566 => x"7487e726",
           567 => x"80d9388a",
           568 => x"13225487",
           569 => x"527387e7",
           570 => x"2680cc38",
           571 => x"810b87c0",
           572 => x"989c0c72",
           573 => x"2287c098",
           574 => x"bc0c8213",
           575 => x"3387c098",
           576 => x"b80c8313",
           577 => x"3387c098",
           578 => x"b40c8413",
           579 => x"3387c098",
           580 => x"b00c8513",
           581 => x"3387c098",
           582 => x"ac0c8613",
           583 => x"3387c098",
           584 => x"a80c7487",
           585 => x"c098a40c",
           586 => x"7387c098",
           587 => x"a00c800b",
           588 => x"87c0989c",
           589 => x"0c805271",
           590 => x"828cec0c",
           591 => x"863d0d04",
           592 => x"f33d0d7f",
           593 => x"5b87c098",
           594 => x"9c5d817d",
           595 => x"0c87c098",
           596 => x"bc085e7d",
           597 => x"7b2387c0",
           598 => x"98b8085a",
           599 => x"79821c34",
           600 => x"87c098b4",
           601 => x"085a7983",
           602 => x"1c3487c0",
           603 => x"98b0085a",
           604 => x"79841c34",
           605 => x"87c098ac",
           606 => x"085a7985",
           607 => x"1c3487c0",
           608 => x"98a8085a",
           609 => x"79861c34",
           610 => x"87c098a4",
           611 => x"085c7b88",
           612 => x"1c2387c0",
           613 => x"98a0085a",
           614 => x"798a1c23",
           615 => x"807d0c79",
           616 => x"83ffff06",
           617 => x"597b83ff",
           618 => x"ff065886",
           619 => x"1b335785",
           620 => x"1b335684",
           621 => x"1b335583",
           622 => x"1b335482",
           623 => x"1b33537d",
           624 => x"83ffff06",
           625 => x"5281f5ec",
           626 => x"5194c93f",
           627 => x"8f3d0d04",
           628 => x"ff3d0d02",
           629 => x"8f053370",
           630 => x"30709f2a",
           631 => x"51525270",
           632 => x"0b0b8289",
           633 => x"9434833d",
           634 => x"0d04fb3d",
           635 => x"0d770b0b",
           636 => x"82899433",
           637 => x"7081ff06",
           638 => x"57555687",
           639 => x"c0948451",
           640 => x"74802e86",
           641 => x"3887c094",
           642 => x"94517008",
           643 => x"70962a70",
           644 => x"81065354",
           645 => x"5270802e",
           646 => x"8c387191",
           647 => x"2a708106",
           648 => x"515170d7",
           649 => x"38728132",
           650 => x"70810651",
           651 => x"5170802e",
           652 => x"8d387193",
           653 => x"2a708106",
           654 => x"515170ff",
           655 => x"be387381",
           656 => x"ff065187",
           657 => x"c0948052",
           658 => x"70802e86",
           659 => x"3887c094",
           660 => x"90527572",
           661 => x"0c75828c",
           662 => x"ec0c873d",
           663 => x"0d04fb3d",
           664 => x"0d029f05",
           665 => x"330b0b82",
           666 => x"89943370",
           667 => x"81ff0657",
           668 => x"555687c0",
           669 => x"94845174",
           670 => x"802e8638",
           671 => x"87c09494",
           672 => x"51700870",
           673 => x"962a7081",
           674 => x"06535452",
           675 => x"70802e8c",
           676 => x"3871912a",
           677 => x"70810651",
           678 => x"5170d738",
           679 => x"72813270",
           680 => x"81065151",
           681 => x"70802e8d",
           682 => x"3871932a",
           683 => x"70810651",
           684 => x"5170ffbe",
           685 => x"387381ff",
           686 => x"065187c0",
           687 => x"94805270",
           688 => x"802e8638",
           689 => x"87c09490",
           690 => x"5275720c",
           691 => x"873d0d04",
           692 => x"f93d0d79",
           693 => x"54807433",
           694 => x"7081ff06",
           695 => x"53535770",
           696 => x"772e80fe",
           697 => x"387181ff",
           698 => x"0681150b",
           699 => x"0b828994",
           700 => x"337081ff",
           701 => x"06595755",
           702 => x"5887c094",
           703 => x"84517580",
           704 => x"2e863887",
           705 => x"c0949451",
           706 => x"70087096",
           707 => x"2a708106",
           708 => x"53545270",
           709 => x"802e8c38",
           710 => x"71912a70",
           711 => x"81065151",
           712 => x"70d73872",
           713 => x"81327081",
           714 => x"06515170",
           715 => x"802e8d38",
           716 => x"71932a70",
           717 => x"81065151",
           718 => x"70ffbe38",
           719 => x"7481ff06",
           720 => x"5187c094",
           721 => x"80527080",
           722 => x"2e863887",
           723 => x"c0949052",
           724 => x"77720c81",
           725 => x"17743370",
           726 => x"81ff0653",
           727 => x"535770ff",
           728 => x"84387682",
           729 => x"8cec0c89",
           730 => x"3d0d04fe",
           731 => x"3d0d0b0b",
           732 => x"82899433",
           733 => x"7081ff06",
           734 => x"545287c0",
           735 => x"94845172",
           736 => x"802e8638",
           737 => x"87c09494",
           738 => x"51700870",
           739 => x"822a7081",
           740 => x"06515151",
           741 => x"70802ee2",
           742 => x"387181ff",
           743 => x"065187c0",
           744 => x"94805270",
           745 => x"802e8638",
           746 => x"87c09490",
           747 => x"52710870",
           748 => x"81ff0682",
           749 => x"8cec0c51",
           750 => x"843d0d04",
           751 => x"fe3d0d0b",
           752 => x"0b828994",
           753 => x"337081ff",
           754 => x"06525387",
           755 => x"c0948452",
           756 => x"70802e86",
           757 => x"3887c094",
           758 => x"94527108",
           759 => x"70822a70",
           760 => x"81065151",
           761 => x"51ff5270",
           762 => x"802ea038",
           763 => x"7281ff06",
           764 => x"5187c094",
           765 => x"80527080",
           766 => x"2e863887",
           767 => x"c0949052",
           768 => x"71087098",
           769 => x"2b70982c",
           770 => x"51535171",
           771 => x"828cec0c",
           772 => x"843d0d04",
           773 => x"ff3d0d87",
           774 => x"c09e8008",
           775 => x"709c2a8a",
           776 => x"06515170",
           777 => x"802e84b4",
           778 => x"3887c09e",
           779 => x"a4088289",
           780 => x"980c87c0",
           781 => x"9ea80882",
           782 => x"899c0c87",
           783 => x"c09e9408",
           784 => x"8289a00c",
           785 => x"87c09e98",
           786 => x"088289a4",
           787 => x"0c87c09e",
           788 => x"9c088289",
           789 => x"a80c87c0",
           790 => x"9ea00882",
           791 => x"89ac0c87",
           792 => x"c09eac08",
           793 => x"8289b00c",
           794 => x"87c09eb0",
           795 => x"088289b4",
           796 => x"0c87c09e",
           797 => x"b4088289",
           798 => x"b80c87c0",
           799 => x"9eb80882",
           800 => x"89bc0c87",
           801 => x"c09ebc08",
           802 => x"8289c00c",
           803 => x"87c09ec0",
           804 => x"088289c4",
           805 => x"0c87c09e",
           806 => x"c4088289",
           807 => x"c80c87c0",
           808 => x"9e800851",
           809 => x"708289cc",
           810 => x"2387c09e",
           811 => x"84088289",
           812 => x"d00c87c0",
           813 => x"9e880882",
           814 => x"89d40c87",
           815 => x"c09e8c08",
           816 => x"8289d80c",
           817 => x"810b8289",
           818 => x"dc34800b",
           819 => x"87c09e90",
           820 => x"08708480",
           821 => x"0a065152",
           822 => x"5270802e",
           823 => x"83388152",
           824 => x"718289dd",
           825 => x"34800b87",
           826 => x"c09e9008",
           827 => x"7088800a",
           828 => x"06515252",
           829 => x"70802e83",
           830 => x"38815271",
           831 => x"8289de34",
           832 => x"800b87c0",
           833 => x"9e900870",
           834 => x"90800a06",
           835 => x"51525270",
           836 => x"802e8338",
           837 => x"81527182",
           838 => x"89df3480",
           839 => x"0b87c09e",
           840 => x"90087088",
           841 => x"80800651",
           842 => x"52527080",
           843 => x"2e833881",
           844 => x"52718289",
           845 => x"e034800b",
           846 => x"87c09e90",
           847 => x"0870a080",
           848 => x"80065152",
           849 => x"5270802e",
           850 => x"83388152",
           851 => x"718289e1",
           852 => x"34800b87",
           853 => x"c09e9008",
           854 => x"70908080",
           855 => x"06515252",
           856 => x"70802e83",
           857 => x"38815271",
           858 => x"8289e234",
           859 => x"800b87c0",
           860 => x"9e900870",
           861 => x"84808006",
           862 => x"51525270",
           863 => x"802e8338",
           864 => x"81527182",
           865 => x"89e33480",
           866 => x"0b87c09e",
           867 => x"90087082",
           868 => x"80800651",
           869 => x"52527080",
           870 => x"2e833881",
           871 => x"52718289",
           872 => x"e434800b",
           873 => x"87c09e90",
           874 => x"08708180",
           875 => x"80065152",
           876 => x"5270802e",
           877 => x"83388152",
           878 => x"718289e5",
           879 => x"34800b87",
           880 => x"c09e9008",
           881 => x"7080c080",
           882 => x"06515252",
           883 => x"70802e83",
           884 => x"38815271",
           885 => x"8289e634",
           886 => x"800b87c0",
           887 => x"9e900870",
           888 => x"a0800651",
           889 => x"52527080",
           890 => x"2e833881",
           891 => x"52718289",
           892 => x"e73487c0",
           893 => x"9e900870",
           894 => x"98800670",
           895 => x"8a2a5151",
           896 => x"51708289",
           897 => x"e834800b",
           898 => x"87c09e90",
           899 => x"08708480",
           900 => x"06515252",
           901 => x"70802e83",
           902 => x"38815271",
           903 => x"8289e934",
           904 => x"87c09e90",
           905 => x"087083f0",
           906 => x"0670842a",
           907 => x"51515170",
           908 => x"8289ea34",
           909 => x"800b87c0",
           910 => x"9e900870",
           911 => x"88065152",
           912 => x"5270802e",
           913 => x"83388152",
           914 => x"718289eb",
           915 => x"3487c09e",
           916 => x"90087087",
           917 => x"06515170",
           918 => x"8289ec34",
           919 => x"833d0d04",
           920 => x"fb3d0d81",
           921 => x"f6845185",
           922 => x"c73f8289",
           923 => x"dc335473",
           924 => x"802e8838",
           925 => x"81f69851",
           926 => x"85b63f81",
           927 => x"f6ac5185",
           928 => x"af3f8289",
           929 => x"de335473",
           930 => x"802e9338",
           931 => x"8289b808",
           932 => x"8289bc08",
           933 => x"11545281",
           934 => x"f6c4518a",
           935 => x"f73f8289",
           936 => x"e3335473",
           937 => x"802e9338",
           938 => x"8289b008",
           939 => x"8289b408",
           940 => x"11545281",
           941 => x"f6e0518a",
           942 => x"db3f8289",
           943 => x"e0335473",
           944 => x"802e9338",
           945 => x"82899808",
           946 => x"82899c08",
           947 => x"11545281",
           948 => x"f6fc518a",
           949 => x"bf3f8289",
           950 => x"e1335473",
           951 => x"802e9338",
           952 => x"8289a008",
           953 => x"8289a408",
           954 => x"11545281",
           955 => x"f798518a",
           956 => x"a33f8289",
           957 => x"e2335473",
           958 => x"802e9338",
           959 => x"8289a808",
           960 => x"8289ac08",
           961 => x"11545281",
           962 => x"f7b4518a",
           963 => x"873f8289",
           964 => x"e7335473",
           965 => x"802e8d38",
           966 => x"8289e833",
           967 => x"5281f7d0",
           968 => x"5189f13f",
           969 => x"8289eb33",
           970 => x"5473802e",
           971 => x"8d388289",
           972 => x"ec335281",
           973 => x"f7f05189",
           974 => x"db3f8289",
           975 => x"e9335473",
           976 => x"802e8d38",
           977 => x"8289ea33",
           978 => x"5281f890",
           979 => x"5189c53f",
           980 => x"8289dd33",
           981 => x"5473802e",
           982 => x"883881f8",
           983 => x"b05183d0",
           984 => x"3f8289df",
           985 => x"33547380",
           986 => x"2e883881",
           987 => x"f8c45183",
           988 => x"bf3f8289",
           989 => x"e4335473",
           990 => x"802e8838",
           991 => x"81f8d051",
           992 => x"83ae3f82",
           993 => x"89e53354",
           994 => x"73802e88",
           995 => x"3881f8dc",
           996 => x"51839d3f",
           997 => x"8289e633",
           998 => x"5473802e",
           999 => x"883881f8",
          1000 => x"e851838c",
          1001 => x"3f81f8f4",
          1002 => x"5183853f",
          1003 => x"8289c008",
          1004 => x"5281f980",
          1005 => x"5188dd3f",
          1006 => x"8289c408",
          1007 => x"5281f9a8",
          1008 => x"5188d13f",
          1009 => x"8289c808",
          1010 => x"5281f9d0",
          1011 => x"5188c53f",
          1012 => x"81f9f851",
          1013 => x"82da3f82",
          1014 => x"89cc2252",
          1015 => x"81fa8051",
          1016 => x"88b23f82",
          1017 => x"89d00856",
          1018 => x"bd84c052",
          1019 => x"7551eac6",
          1020 => x"3f828cec",
          1021 => x"08bd84c0",
          1022 => x"29767131",
          1023 => x"5454828c",
          1024 => x"ec085281",
          1025 => x"faa85188",
          1026 => x"8b3f8289",
          1027 => x"e3335473",
          1028 => x"802ea838",
          1029 => x"8289d408",
          1030 => x"56bd84c0",
          1031 => x"527551ea",
          1032 => x"953f828c",
          1033 => x"ec08bd84",
          1034 => x"c0297671",
          1035 => x"31545482",
          1036 => x"8cec0852",
          1037 => x"81fad451",
          1038 => x"87da3f82",
          1039 => x"89de3354",
          1040 => x"73802ea8",
          1041 => x"388289d8",
          1042 => x"0856bd84",
          1043 => x"c0527551",
          1044 => x"e9e43f82",
          1045 => x"8cec08bd",
          1046 => x"84c02976",
          1047 => x"71315454",
          1048 => x"828cec08",
          1049 => x"5281fb80",
          1050 => x"5187a93f",
          1051 => x"8286e451",
          1052 => x"81be3f87",
          1053 => x"3d0d04fe",
          1054 => x"3d0d0292",
          1055 => x"0533ff05",
          1056 => x"52718426",
          1057 => x"ac387184",
          1058 => x"290b0b81",
          1059 => x"f5880552",
          1060 => x"71080481",
          1061 => x"fbac519d",
          1062 => x"3981fbb4",
          1063 => x"51973981",
          1064 => x"fbbc5191",
          1065 => x"3981fbc4",
          1066 => x"518b3981",
          1067 => x"fbc85185",
          1068 => x"3981fbd0",
          1069 => x"5180f93f",
          1070 => x"843d0d04",
          1071 => x"7188800c",
          1072 => x"04800b87",
          1073 => x"c096840c",
          1074 => x"048289f0",
          1075 => x"0887c096",
          1076 => x"840c04fe",
          1077 => x"3d0d0293",
          1078 => x"05335372",
          1079 => x"8a2e0981",
          1080 => x"0685388d",
          1081 => x"51ed3f82",
          1082 => x"8d840852",
          1083 => x"71802e90",
          1084 => x"38727234",
          1085 => x"828d8408",
          1086 => x"8105828d",
          1087 => x"840c8f39",
          1088 => x"828cfc08",
          1089 => x"5271802e",
          1090 => x"85387251",
          1091 => x"712d843d",
          1092 => x"0d04fe3d",
          1093 => x"0d029705",
          1094 => x"33828cfc",
          1095 => x"0876828c",
          1096 => x"fc0c5451",
          1097 => x"ffad3f72",
          1098 => x"828cfc0c",
          1099 => x"843d0d04",
          1100 => x"fd3d0d75",
          1101 => x"54733370",
          1102 => x"81ff0653",
          1103 => x"5371802e",
          1104 => x"8e387281",
          1105 => x"ff065181",
          1106 => x"1454ff87",
          1107 => x"3fe73985",
          1108 => x"3d0d04fc",
          1109 => x"3d0d7782",
          1110 => x"8cfc0878",
          1111 => x"828cfc0c",
          1112 => x"56547333",
          1113 => x"7081ff06",
          1114 => x"53537180",
          1115 => x"2e8e3872",
          1116 => x"81ff0651",
          1117 => x"811454fe",
          1118 => x"da3fe739",
          1119 => x"74828cfc",
          1120 => x"0c863d0d",
          1121 => x"04ec3d0d",
          1122 => x"66685959",
          1123 => x"78708105",
          1124 => x"5a335675",
          1125 => x"802e84f8",
          1126 => x"3875a52e",
          1127 => x"09810682",
          1128 => x"de388070",
          1129 => x"7a708105",
          1130 => x"5c33585b",
          1131 => x"5b75b02e",
          1132 => x"09810685",
          1133 => x"38815a8b",
          1134 => x"3975ad2e",
          1135 => x"0981068a",
          1136 => x"38825a78",
          1137 => x"7081055a",
          1138 => x"335675aa",
          1139 => x"2e098106",
          1140 => x"92387784",
          1141 => x"1971087b",
          1142 => x"7081055d",
          1143 => x"33595d59",
          1144 => x"539d39d0",
          1145 => x"16537289",
          1146 => x"2695387a",
          1147 => x"88297b10",
          1148 => x"057605d0",
          1149 => x"05797081",
          1150 => x"055b3357",
          1151 => x"5be53975",
          1152 => x"80ec3270",
          1153 => x"30707207",
          1154 => x"80257880",
          1155 => x"cc327030",
          1156 => x"70720780",
          1157 => x"25730753",
          1158 => x"54585155",
          1159 => x"5373802e",
          1160 => x"8c387984",
          1161 => x"07797081",
          1162 => x"055b3357",
          1163 => x"5a75802e",
          1164 => x"83de3875",
          1165 => x"5480e076",
          1166 => x"278938e0",
          1167 => x"167081ff",
          1168 => x"06555373",
          1169 => x"80cf2e81",
          1170 => x"aa387380",
          1171 => x"cf24a238",
          1172 => x"7380c32e",
          1173 => x"818e3873",
          1174 => x"80c3248b",
          1175 => x"387380c2",
          1176 => x"2e818c38",
          1177 => x"81993973",
          1178 => x"80c42e81",
          1179 => x"8a38818f",
          1180 => x"397380d5",
          1181 => x"2e818038",
          1182 => x"7380d524",
          1183 => x"8a387380",
          1184 => x"d32e8e38",
          1185 => x"80f93973",
          1186 => x"80d82e80",
          1187 => x"ee3880ef",
          1188 => x"39778419",
          1189 => x"71085659",
          1190 => x"53807433",
          1191 => x"54557275",
          1192 => x"2e8d3881",
          1193 => x"15701570",
          1194 => x"33515455",
          1195 => x"72f53879",
          1196 => x"812a5690",
          1197 => x"39748116",
          1198 => x"5653727b",
          1199 => x"278f38a0",
          1200 => x"51fc903f",
          1201 => x"75810653",
          1202 => x"72802ee9",
          1203 => x"387351fc",
          1204 => x"df3f7481",
          1205 => x"16565372",
          1206 => x"7b27fdb0",
          1207 => x"38a051fb",
          1208 => x"f23fef39",
          1209 => x"77841983",
          1210 => x"12335359",
          1211 => x"53933982",
          1212 => x"5c953988",
          1213 => x"5c91398a",
          1214 => x"5c8d3990",
          1215 => x"5c893975",
          1216 => x"51fbd03f",
          1217 => x"fd863979",
          1218 => x"822a7081",
          1219 => x"06515372",
          1220 => x"802e8838",
          1221 => x"77841959",
          1222 => x"53863984",
          1223 => x"18785458",
          1224 => x"72087480",
          1225 => x"c4327030",
          1226 => x"70720780",
          1227 => x"25515555",
          1228 => x"55748025",
          1229 => x"8d387280",
          1230 => x"2e883874",
          1231 => x"307a9007",
          1232 => x"5b55800b",
          1233 => x"8f3d5e57",
          1234 => x"7b527451",
          1235 => x"e49b3f82",
          1236 => x"8cec0881",
          1237 => x"ff067c53",
          1238 => x"755254e3",
          1239 => x"d93f828c",
          1240 => x"ec085589",
          1241 => x"74279238",
          1242 => x"a7145375",
          1243 => x"80f82e84",
          1244 => x"38871453",
          1245 => x"7281ff06",
          1246 => x"54b01453",
          1247 => x"727d7081",
          1248 => x"055f3481",
          1249 => x"17753070",
          1250 => x"77079f2a",
          1251 => x"51545776",
          1252 => x"9f268538",
          1253 => x"72ffb138",
          1254 => x"79842a70",
          1255 => x"81065153",
          1256 => x"72802e8e",
          1257 => x"38963d77",
          1258 => x"05e00553",
          1259 => x"ad733481",
          1260 => x"1757767a",
          1261 => x"81065455",
          1262 => x"b0547283",
          1263 => x"38a05479",
          1264 => x"812a7081",
          1265 => x"06545672",
          1266 => x"9f388117",
          1267 => x"55767b27",
          1268 => x"97387351",
          1269 => x"f9fd3f75",
          1270 => x"81065372",
          1271 => x"8b387481",
          1272 => x"1656537a",
          1273 => x"7326eb38",
          1274 => x"963d7705",
          1275 => x"e00553ff",
          1276 => x"17ff1470",
          1277 => x"33535457",
          1278 => x"f9d93f76",
          1279 => x"f2387481",
          1280 => x"16565372",
          1281 => x"7b27fb84",
          1282 => x"38a051f9",
          1283 => x"c63fef39",
          1284 => x"963d0d04",
          1285 => x"fd3d0d86",
          1286 => x"3d707084",
          1287 => x"05520855",
          1288 => x"527351fa",
          1289 => x"e03f853d",
          1290 => x"0d04fe3d",
          1291 => x"0d74828d",
          1292 => x"840c853d",
          1293 => x"88055275",
          1294 => x"51faca3f",
          1295 => x"828d8408",
          1296 => x"53807334",
          1297 => x"800b828d",
          1298 => x"840c843d",
          1299 => x"0d04fd3d",
          1300 => x"0d828cfc",
          1301 => x"0876828c",
          1302 => x"fc0c873d",
          1303 => x"88055377",
          1304 => x"5253faa1",
          1305 => x"3f72828c",
          1306 => x"fc0c853d",
          1307 => x"0d04fb3d",
          1308 => x"0d777982",
          1309 => x"8d800870",
          1310 => x"56545755",
          1311 => x"80547180",
          1312 => x"2e80e038",
          1313 => x"828d8008",
          1314 => x"52712d82",
          1315 => x"8cec0881",
          1316 => x"ff065372",
          1317 => x"802e80cb",
          1318 => x"38728d2e",
          1319 => x"b9387288",
          1320 => x"32703070",
          1321 => x"80255151",
          1322 => x"5273802e",
          1323 => x"8b387180",
          1324 => x"2e8638ff",
          1325 => x"14549739",
          1326 => x"9f7325c8",
          1327 => x"38ff1652",
          1328 => x"737225c0",
          1329 => x"38741452",
          1330 => x"72723481",
          1331 => x"14547251",
          1332 => x"f8813fff",
          1333 => x"af397315",
          1334 => x"52807234",
          1335 => x"8a51f7f3",
          1336 => x"3f815372",
          1337 => x"828cec0c",
          1338 => x"873d0d04",
          1339 => x"fe3d0d82",
          1340 => x"8d800875",
          1341 => x"828d800c",
          1342 => x"77537652",
          1343 => x"53feef3f",
          1344 => x"72828d80",
          1345 => x"0c843d0d",
          1346 => x"04f83d0d",
          1347 => x"7a7c5a56",
          1348 => x"80707a0c",
          1349 => x"58750870",
          1350 => x"33555373",
          1351 => x"a02e0981",
          1352 => x"06873881",
          1353 => x"13760ced",
          1354 => x"3973ad2e",
          1355 => x"0981068e",
          1356 => x"38817608",
          1357 => x"11770c76",
          1358 => x"08703356",
          1359 => x"545873b0",
          1360 => x"2e098106",
          1361 => x"80c23875",
          1362 => x"08810576",
          1363 => x"0c750870",
          1364 => x"33555373",
          1365 => x"80e22e8b",
          1366 => x"38905773",
          1367 => x"80f82e85",
          1368 => x"388f3982",
          1369 => x"57811376",
          1370 => x"0c750870",
          1371 => x"335553ac",
          1372 => x"398155a0",
          1373 => x"742780fa",
          1374 => x"38d01453",
          1375 => x"80558857",
          1376 => x"89732798",
          1377 => x"3880eb39",
          1378 => x"d0145380",
          1379 => x"55728926",
          1380 => x"80e03886",
          1381 => x"39805580",
          1382 => x"d9398a57",
          1383 => x"8055a074",
          1384 => x"2780c238",
          1385 => x"80e07427",
          1386 => x"8938e014",
          1387 => x"7081ff06",
          1388 => x"5553d014",
          1389 => x"7081ff06",
          1390 => x"55539074",
          1391 => x"278e38f9",
          1392 => x"147081ff",
          1393 => x"06555389",
          1394 => x"7427ca38",
          1395 => x"737727c5",
          1396 => x"38747729",
          1397 => x"14760881",
          1398 => x"05770c76",
          1399 => x"08703356",
          1400 => x"5455ffba",
          1401 => x"3977802e",
          1402 => x"84387430",
          1403 => x"5574790c",
          1404 => x"81557482",
          1405 => x"8cec0c8a",
          1406 => x"3d0d04f8",
          1407 => x"3d0d7a7c",
          1408 => x"5a568070",
          1409 => x"7a0c5875",
          1410 => x"08703355",
          1411 => x"5373a02e",
          1412 => x"09810687",
          1413 => x"38811376",
          1414 => x"0ced3973",
          1415 => x"ad2e0981",
          1416 => x"068e3881",
          1417 => x"76081177",
          1418 => x"0c760870",
          1419 => x"33565458",
          1420 => x"73b02e09",
          1421 => x"810680c2",
          1422 => x"38750881",
          1423 => x"05760c75",
          1424 => x"08703355",
          1425 => x"537380e2",
          1426 => x"2e8b3890",
          1427 => x"577380f8",
          1428 => x"2e85388f",
          1429 => x"39825781",
          1430 => x"13760c75",
          1431 => x"08703355",
          1432 => x"53ac3981",
          1433 => x"55a07427",
          1434 => x"80fa38d0",
          1435 => x"14538055",
          1436 => x"88578973",
          1437 => x"27983880",
          1438 => x"eb39d014",
          1439 => x"53805572",
          1440 => x"892680e0",
          1441 => x"38863980",
          1442 => x"5580d939",
          1443 => x"8a578055",
          1444 => x"a0742780",
          1445 => x"c23880e0",
          1446 => x"74278938",
          1447 => x"e0147081",
          1448 => x"ff065553",
          1449 => x"d0147081",
          1450 => x"ff065553",
          1451 => x"9074278e",
          1452 => x"38f91470",
          1453 => x"81ff0655",
          1454 => x"53897427",
          1455 => x"ca387377",
          1456 => x"27c53874",
          1457 => x"77291476",
          1458 => x"08810577",
          1459 => x"0c760870",
          1460 => x"33565455",
          1461 => x"ffba3977",
          1462 => x"802e8438",
          1463 => x"74305574",
          1464 => x"790c8155",
          1465 => x"74828cec",
          1466 => x"0c8a3d0d",
          1467 => x"04ff3d0d",
          1468 => x"028f0533",
          1469 => x"51815270",
          1470 => x"72268738",
          1471 => x"8289f411",
          1472 => x"33527182",
          1473 => x"8cec0c83",
          1474 => x"3d0d04fc",
          1475 => x"3d0d029b",
          1476 => x"05330284",
          1477 => x"059f0533",
          1478 => x"56538351",
          1479 => x"72812680",
          1480 => x"e0387284",
          1481 => x"2b87c092",
          1482 => x"8c115351",
          1483 => x"88547480",
          1484 => x"2e843881",
          1485 => x"88547372",
          1486 => x"0c87c092",
          1487 => x"8c115181",
          1488 => x"710c850b",
          1489 => x"87c0988c",
          1490 => x"0c705271",
          1491 => x"08708206",
          1492 => x"51517080",
          1493 => x"2e8a3887",
          1494 => x"c0988c08",
          1495 => x"5170ec38",
          1496 => x"7108fc80",
          1497 => x"80065271",
          1498 => x"923887c0",
          1499 => x"988c0851",
          1500 => x"70802e87",
          1501 => x"38718289",
          1502 => x"f4143482",
          1503 => x"89f41333",
          1504 => x"5170828c",
          1505 => x"ec0c863d",
          1506 => x"0d04f33d",
          1507 => x"0d606264",
          1508 => x"028c05bf",
          1509 => x"05335740",
          1510 => x"585b8374",
          1511 => x"525afecd",
          1512 => x"3f828cec",
          1513 => x"0881067a",
          1514 => x"54527181",
          1515 => x"be387172",
          1516 => x"75842b87",
          1517 => x"c0928011",
          1518 => x"87c0928c",
          1519 => x"1287c092",
          1520 => x"8413415a",
          1521 => x"40575a58",
          1522 => x"850b87c0",
          1523 => x"988c0c76",
          1524 => x"7d0c8476",
          1525 => x"0c750870",
          1526 => x"852a7081",
          1527 => x"06515354",
          1528 => x"71802e8e",
          1529 => x"387b0852",
          1530 => x"717b7081",
          1531 => x"055d3481",
          1532 => x"19598074",
          1533 => x"a2065353",
          1534 => x"71732e83",
          1535 => x"38815378",
          1536 => x"83ff268f",
          1537 => x"3872802e",
          1538 => x"8a3887c0",
          1539 => x"988c0852",
          1540 => x"71c33887",
          1541 => x"c0988c08",
          1542 => x"5271802e",
          1543 => x"87387884",
          1544 => x"802e9938",
          1545 => x"81760c87",
          1546 => x"c0928c15",
          1547 => x"53720870",
          1548 => x"82065152",
          1549 => x"71f738ff",
          1550 => x"1a5a8d39",
          1551 => x"84801781",
          1552 => x"197081ff",
          1553 => x"065a5357",
          1554 => x"79802e90",
          1555 => x"3873fc80",
          1556 => x"80065271",
          1557 => x"87387d78",
          1558 => x"26feed38",
          1559 => x"73fc8080",
          1560 => x"06527180",
          1561 => x"2e833881",
          1562 => x"52715372",
          1563 => x"828cec0c",
          1564 => x"8f3d0d04",
          1565 => x"f33d0d60",
          1566 => x"6264028c",
          1567 => x"05bf0533",
          1568 => x"5740585b",
          1569 => x"83598074",
          1570 => x"5258fce1",
          1571 => x"3f828cec",
          1572 => x"08810679",
          1573 => x"54527178",
          1574 => x"2e098106",
          1575 => x"81b13877",
          1576 => x"74842b87",
          1577 => x"c0928011",
          1578 => x"87c0928c",
          1579 => x"1287c092",
          1580 => x"84134059",
          1581 => x"5f565a85",
          1582 => x"0b87c098",
          1583 => x"8c0c767d",
          1584 => x"0c82760c",
          1585 => x"80587508",
          1586 => x"70842a70",
          1587 => x"81065153",
          1588 => x"5471802e",
          1589 => x"8c387a70",
          1590 => x"81055c33",
          1591 => x"7c0c8118",
          1592 => x"5873812a",
          1593 => x"70810651",
          1594 => x"5271802e",
          1595 => x"8a3887c0",
          1596 => x"988c0852",
          1597 => x"71d03887",
          1598 => x"c0988c08",
          1599 => x"5271802e",
          1600 => x"87387784",
          1601 => x"802e9938",
          1602 => x"81760c87",
          1603 => x"c0928c15",
          1604 => x"53720870",
          1605 => x"82065152",
          1606 => x"71f738ff",
          1607 => x"19598d39",
          1608 => x"811a7081",
          1609 => x"ff068480",
          1610 => x"19595b52",
          1611 => x"78802e90",
          1612 => x"3873fc80",
          1613 => x"80065271",
          1614 => x"87387d7a",
          1615 => x"26fef838",
          1616 => x"73fc8080",
          1617 => x"06527180",
          1618 => x"2e833881",
          1619 => x"52715372",
          1620 => x"828cec0c",
          1621 => x"8f3d0d04",
          1622 => x"fa3d0d7a",
          1623 => x"028405a3",
          1624 => x"05330288",
          1625 => x"05a70533",
          1626 => x"71545456",
          1627 => x"57fafe3f",
          1628 => x"828cec08",
          1629 => x"81065383",
          1630 => x"547280fe",
          1631 => x"38850b87",
          1632 => x"c0988c0c",
          1633 => x"81567176",
          1634 => x"2e80dc38",
          1635 => x"71762493",
          1636 => x"3874842b",
          1637 => x"87c0928c",
          1638 => x"11545471",
          1639 => x"802e8d38",
          1640 => x"80d43971",
          1641 => x"832e80c6",
          1642 => x"3880cb39",
          1643 => x"72087081",
          1644 => x"2a708106",
          1645 => x"51515271",
          1646 => x"802e8a38",
          1647 => x"87c0988c",
          1648 => x"085271e8",
          1649 => x"3887c098",
          1650 => x"8c085271",
          1651 => x"96388173",
          1652 => x"0c87c092",
          1653 => x"8c145372",
          1654 => x"08708206",
          1655 => x"515271f7",
          1656 => x"38963980",
          1657 => x"56923988",
          1658 => x"800a770c",
          1659 => x"85398180",
          1660 => x"770c7256",
          1661 => x"83398456",
          1662 => x"75547382",
          1663 => x"8cec0c88",
          1664 => x"3d0d04fe",
          1665 => x"3d0d7481",
          1666 => x"11337133",
          1667 => x"71882b07",
          1668 => x"828cec0c",
          1669 => x"5351843d",
          1670 => x"0d04fd3d",
          1671 => x"0d758311",
          1672 => x"33821233",
          1673 => x"71902b71",
          1674 => x"882b0781",
          1675 => x"14337072",
          1676 => x"07882b75",
          1677 => x"33710782",
          1678 => x"8cec0c52",
          1679 => x"53545654",
          1680 => x"52853d0d",
          1681 => x"04ff3d0d",
          1682 => x"73028405",
          1683 => x"92052252",
          1684 => x"52707270",
          1685 => x"81055434",
          1686 => x"70882a51",
          1687 => x"70723483",
          1688 => x"3d0d04ff",
          1689 => x"3d0d7375",
          1690 => x"52527072",
          1691 => x"70810554",
          1692 => x"3470882a",
          1693 => x"51707270",
          1694 => x"81055434",
          1695 => x"70882a51",
          1696 => x"70727081",
          1697 => x"05543470",
          1698 => x"882a5170",
          1699 => x"7234833d",
          1700 => x"0d04fe3d",
          1701 => x"0d767577",
          1702 => x"54545170",
          1703 => x"802e9238",
          1704 => x"71708105",
          1705 => x"53337370",
          1706 => x"81055534",
          1707 => x"ff1151eb",
          1708 => x"39843d0d",
          1709 => x"04fe3d0d",
          1710 => x"75777654",
          1711 => x"52537272",
          1712 => x"70810554",
          1713 => x"34ff1151",
          1714 => x"70f43884",
          1715 => x"3d0d04fc",
          1716 => x"3d0d7877",
          1717 => x"79565653",
          1718 => x"74708105",
          1719 => x"56337470",
          1720 => x"81055633",
          1721 => x"717131ff",
          1722 => x"16565252",
          1723 => x"5272802e",
          1724 => x"86387180",
          1725 => x"2ee23871",
          1726 => x"828cec0c",
          1727 => x"863d0d04",
          1728 => x"fe3d0d74",
          1729 => x"76545189",
          1730 => x"3971732e",
          1731 => x"8a388111",
          1732 => x"51703352",
          1733 => x"71f33870",
          1734 => x"33828cec",
          1735 => x"0c843d0d",
          1736 => x"04800b82",
          1737 => x"8cec0c04",
          1738 => x"800b828c",
          1739 => x"ec0c04f7",
          1740 => x"3d0d7b56",
          1741 => x"800b8317",
          1742 => x"33565a74",
          1743 => x"7a2e80d6",
          1744 => x"388154b0",
          1745 => x"160853b4",
          1746 => x"16705381",
          1747 => x"17335259",
          1748 => x"faa23f82",
          1749 => x"8cec087a",
          1750 => x"2e098106",
          1751 => x"b738828c",
          1752 => x"ec088317",
          1753 => x"34b01608",
          1754 => x"70a41808",
          1755 => x"319c1808",
          1756 => x"59565874",
          1757 => x"77279f38",
          1758 => x"82163355",
          1759 => x"74822e09",
          1760 => x"81069338",
          1761 => x"81547618",
          1762 => x"53785281",
          1763 => x"163351f9",
          1764 => x"e33f8339",
          1765 => x"815a7982",
          1766 => x"8cec0c8b",
          1767 => x"3d0d04fa",
          1768 => x"3d0d787a",
          1769 => x"56568057",
          1770 => x"74b01708",
          1771 => x"2eaf3875",
          1772 => x"51fefc3f",
          1773 => x"828cec08",
          1774 => x"57828cec",
          1775 => x"089f3881",
          1776 => x"547453b4",
          1777 => x"16528116",
          1778 => x"3351f7be",
          1779 => x"3f828cec",
          1780 => x"08802e85",
          1781 => x"38ff5581",
          1782 => x"5774b017",
          1783 => x"0c76828c",
          1784 => x"ec0c883d",
          1785 => x"0d04f83d",
          1786 => x"0d7a7052",
          1787 => x"57fec03f",
          1788 => x"828cec08",
          1789 => x"58828cec",
          1790 => x"08819138",
          1791 => x"76335574",
          1792 => x"832e0981",
          1793 => x"0680f038",
          1794 => x"84173359",
          1795 => x"78812e09",
          1796 => x"810680e3",
          1797 => x"38848053",
          1798 => x"828cec08",
          1799 => x"52b41770",
          1800 => x"5256fd91",
          1801 => x"3f82d4d5",
          1802 => x"5284b217",
          1803 => x"51fc963f",
          1804 => x"848b85a4",
          1805 => x"d2527551",
          1806 => x"fca93f86",
          1807 => x"8a85e4f2",
          1808 => x"52849817",
          1809 => x"51fc9c3f",
          1810 => x"90170852",
          1811 => x"849c1751",
          1812 => x"fc913f8c",
          1813 => x"17085284",
          1814 => x"a01751fc",
          1815 => x"863fa017",
          1816 => x"08810570",
          1817 => x"b0190c79",
          1818 => x"55537552",
          1819 => x"81173351",
          1820 => x"f8823f77",
          1821 => x"84183480",
          1822 => x"53805281",
          1823 => x"173351f9",
          1824 => x"d73f828c",
          1825 => x"ec08802e",
          1826 => x"83388158",
          1827 => x"77828cec",
          1828 => x"0c8a3d0d",
          1829 => x"04fb3d0d",
          1830 => x"77fe1a98",
          1831 => x"1208fe05",
          1832 => x"55565480",
          1833 => x"56747327",
          1834 => x"8d388a14",
          1835 => x"22757129",
          1836 => x"ac160805",
          1837 => x"57537582",
          1838 => x"8cec0c87",
          1839 => x"3d0d04f9",
          1840 => x"3d0d7a7a",
          1841 => x"70085654",
          1842 => x"57817727",
          1843 => x"81df3876",
          1844 => x"98150827",
          1845 => x"81d738ff",
          1846 => x"74335458",
          1847 => x"72822e80",
          1848 => x"f5387282",
          1849 => x"24893872",
          1850 => x"812e8d38",
          1851 => x"81bf3972",
          1852 => x"832e818e",
          1853 => x"3881b639",
          1854 => x"76812a17",
          1855 => x"70892aa4",
          1856 => x"16080553",
          1857 => x"745255fd",
          1858 => x"963f828c",
          1859 => x"ec08819f",
          1860 => x"387483ff",
          1861 => x"0614b411",
          1862 => x"33811770",
          1863 => x"892aa418",
          1864 => x"08055576",
          1865 => x"54575753",
          1866 => x"fcf53f82",
          1867 => x"8cec0880",
          1868 => x"fe387483",
          1869 => x"ff0614b4",
          1870 => x"11337088",
          1871 => x"2b780779",
          1872 => x"81067184",
          1873 => x"2a5c5258",
          1874 => x"51537280",
          1875 => x"e238759f",
          1876 => x"ff065880",
          1877 => x"da397688",
          1878 => x"2aa41508",
          1879 => x"05527351",
          1880 => x"fcbd3f82",
          1881 => x"8cec0880",
          1882 => x"c6387610",
          1883 => x"83fe0674",
          1884 => x"05b40551",
          1885 => x"f98d3f82",
          1886 => x"8cec0883",
          1887 => x"ffff0658",
          1888 => x"ae397687",
          1889 => x"2aa41508",
          1890 => x"05527351",
          1891 => x"fc913f82",
          1892 => x"8cec089b",
          1893 => x"3876822b",
          1894 => x"83fc0674",
          1895 => x"05b40551",
          1896 => x"f8f83f82",
          1897 => x"8cec08f0",
          1898 => x"0a065883",
          1899 => x"39815877",
          1900 => x"828cec0c",
          1901 => x"893d0d04",
          1902 => x"f83d0d7a",
          1903 => x"7c7e5a58",
          1904 => x"56825981",
          1905 => x"7727829e",
          1906 => x"38769817",
          1907 => x"08278296",
          1908 => x"38753353",
          1909 => x"72792e81",
          1910 => x"9d387279",
          1911 => x"24893872",
          1912 => x"812e8d38",
          1913 => x"82803972",
          1914 => x"832e81b8",
          1915 => x"3881f739",
          1916 => x"76812a17",
          1917 => x"70892aa4",
          1918 => x"18080553",
          1919 => x"765255fb",
          1920 => x"9e3f828c",
          1921 => x"ec085982",
          1922 => x"8cec0881",
          1923 => x"d9387483",
          1924 => x"ff0616b4",
          1925 => x"05811678",
          1926 => x"81065956",
          1927 => x"54775376",
          1928 => x"802e8f38",
          1929 => x"77842b9f",
          1930 => x"f0067433",
          1931 => x"8f067107",
          1932 => x"51537274",
          1933 => x"34810b83",
          1934 => x"17347489",
          1935 => x"2aa41708",
          1936 => x"05527551",
          1937 => x"fad93f82",
          1938 => x"8cec0859",
          1939 => x"828cec08",
          1940 => x"81943874",
          1941 => x"83ff0616",
          1942 => x"b4057884",
          1943 => x"2a545476",
          1944 => x"8f387788",
          1945 => x"2a743381",
          1946 => x"f006718f",
          1947 => x"06075153",
          1948 => x"72743480",
          1949 => x"ec397688",
          1950 => x"2aa41708",
          1951 => x"05527551",
          1952 => x"fa9d3f82",
          1953 => x"8cec0859",
          1954 => x"828cec08",
          1955 => x"80d83877",
          1956 => x"83ffff06",
          1957 => x"52761083",
          1958 => x"fe067605",
          1959 => x"b40551f7",
          1960 => x"a43fbe39",
          1961 => x"76872aa4",
          1962 => x"17080552",
          1963 => x"7551f9ef",
          1964 => x"3f828cec",
          1965 => x"0859828c",
          1966 => x"ec08ab38",
          1967 => x"77f00a06",
          1968 => x"77822b83",
          1969 => x"fc067018",
          1970 => x"b4057054",
          1971 => x"515454f6",
          1972 => x"c93f828c",
          1973 => x"ec088f0a",
          1974 => x"06740752",
          1975 => x"7251f783",
          1976 => x"3f810b83",
          1977 => x"17347882",
          1978 => x"8cec0c8a",
          1979 => x"3d0d04f8",
          1980 => x"3d0d7a7c",
          1981 => x"7e720859",
          1982 => x"56565981",
          1983 => x"7527a438",
          1984 => x"74981708",
          1985 => x"279d3873",
          1986 => x"802eaa38",
          1987 => x"ff537352",
          1988 => x"7551fda4",
          1989 => x"3f828cec",
          1990 => x"0854828c",
          1991 => x"ec0880f2",
          1992 => x"38933982",
          1993 => x"5480eb39",
          1994 => x"815480e6",
          1995 => x"39828cec",
          1996 => x"085480de",
          1997 => x"39745278",
          1998 => x"51fb843f",
          1999 => x"828cec08",
          2000 => x"58828cec",
          2001 => x"08802e80",
          2002 => x"c738828c",
          2003 => x"ec08812e",
          2004 => x"d238828c",
          2005 => x"ec08ff2e",
          2006 => x"cf388053",
          2007 => x"74527551",
          2008 => x"fcd63f82",
          2009 => x"8cec08c5",
          2010 => x"38981608",
          2011 => x"fe119018",
          2012 => x"08575557",
          2013 => x"74742790",
          2014 => x"38811590",
          2015 => x"170c8416",
          2016 => x"33810754",
          2017 => x"73841734",
          2018 => x"77557678",
          2019 => x"26ffa638",
          2020 => x"80547382",
          2021 => x"8cec0c8a",
          2022 => x"3d0d04f6",
          2023 => x"3d0d7c7e",
          2024 => x"7108595b",
          2025 => x"5b799538",
          2026 => x"8c170858",
          2027 => x"77802e88",
          2028 => x"38981708",
          2029 => x"7826b238",
          2030 => x"8158ae39",
          2031 => x"79527a51",
          2032 => x"f9fd3f81",
          2033 => x"5574828c",
          2034 => x"ec082782",
          2035 => x"e038828c",
          2036 => x"ec085582",
          2037 => x"8cec08ff",
          2038 => x"2e82d238",
          2039 => x"98170882",
          2040 => x"8cec0826",
          2041 => x"82c73879",
          2042 => x"58901708",
          2043 => x"70565473",
          2044 => x"802e82b9",
          2045 => x"38777a2e",
          2046 => x"09810680",
          2047 => x"e238811a",
          2048 => x"56981708",
          2049 => x"76268338",
          2050 => x"82567552",
          2051 => x"7a51f9af",
          2052 => x"3f805982",
          2053 => x"8cec0881",
          2054 => x"2e098106",
          2055 => x"8638828c",
          2056 => x"ec085982",
          2057 => x"8cec0809",
          2058 => x"70307072",
          2059 => x"07802570",
          2060 => x"7c07828c",
          2061 => x"ec085451",
          2062 => x"51555573",
          2063 => x"81ef3882",
          2064 => x"8cec0880",
          2065 => x"2e95388c",
          2066 => x"17085481",
          2067 => x"74279038",
          2068 => x"73981808",
          2069 => x"27893873",
          2070 => x"58853975",
          2071 => x"80db3877",
          2072 => x"56811656",
          2073 => x"98170876",
          2074 => x"26893882",
          2075 => x"56757826",
          2076 => x"81ac3875",
          2077 => x"527a51f8",
          2078 => x"c63f828c",
          2079 => x"ec08802e",
          2080 => x"b8388059",
          2081 => x"828cec08",
          2082 => x"812e0981",
          2083 => x"06863882",
          2084 => x"8cec0859",
          2085 => x"828cec08",
          2086 => x"09703070",
          2087 => x"72078025",
          2088 => x"707c0751",
          2089 => x"51555573",
          2090 => x"80f83875",
          2091 => x"782e0981",
          2092 => x"06ffae38",
          2093 => x"735580f5",
          2094 => x"39ff5375",
          2095 => x"527651f9",
          2096 => x"f73f828c",
          2097 => x"ec08828c",
          2098 => x"ec083070",
          2099 => x"828cec08",
          2100 => x"07802551",
          2101 => x"55557980",
          2102 => x"2e943873",
          2103 => x"802e8f38",
          2104 => x"75537952",
          2105 => x"7651f9d0",
          2106 => x"3f828cec",
          2107 => x"085574a5",
          2108 => x"38758c18",
          2109 => x"0c981708",
          2110 => x"fe059018",
          2111 => x"08565474",
          2112 => x"74268638",
          2113 => x"ff159018",
          2114 => x"0c841733",
          2115 => x"81075473",
          2116 => x"84183497",
          2117 => x"39ff5674",
          2118 => x"812e9038",
          2119 => x"8c398055",
          2120 => x"8c39828c",
          2121 => x"ec085585",
          2122 => x"39815675",
          2123 => x"5574828c",
          2124 => x"ec0c8c3d",
          2125 => x"0d04f83d",
          2126 => x"0d7a7052",
          2127 => x"55f3f03f",
          2128 => x"828cec08",
          2129 => x"58815682",
          2130 => x"8cec0880",
          2131 => x"d8387b52",
          2132 => x"7451f6c1",
          2133 => x"3f828cec",
          2134 => x"08828cec",
          2135 => x"08b0170c",
          2136 => x"59848053",
          2137 => x"7752b415",
          2138 => x"705257f2",
          2139 => x"c83f7756",
          2140 => x"84398116",
          2141 => x"568a1522",
          2142 => x"58757827",
          2143 => x"97388154",
          2144 => x"75195376",
          2145 => x"52811533",
          2146 => x"51ede93f",
          2147 => x"828cec08",
          2148 => x"802edf38",
          2149 => x"8a152276",
          2150 => x"32703070",
          2151 => x"7207709f",
          2152 => x"2a535156",
          2153 => x"5675828c",
          2154 => x"ec0c8a3d",
          2155 => x"0d04f83d",
          2156 => x"0d7a7c71",
          2157 => x"08585657",
          2158 => x"74f0800a",
          2159 => x"2680f138",
          2160 => x"749f0653",
          2161 => x"7280e938",
          2162 => x"7490180c",
          2163 => x"88170854",
          2164 => x"73aa3875",
          2165 => x"33538273",
          2166 => x"278838a8",
          2167 => x"16085473",
          2168 => x"9b387485",
          2169 => x"2a53820b",
          2170 => x"8817225a",
          2171 => x"58727927",
          2172 => x"80fe38a8",
          2173 => x"16089818",
          2174 => x"0c80cd39",
          2175 => x"8a162270",
          2176 => x"892b5458",
          2177 => x"727526b2",
          2178 => x"38735276",
          2179 => x"51f5b03f",
          2180 => x"828cec08",
          2181 => x"54828cec",
          2182 => x"08ff2ebd",
          2183 => x"38810b82",
          2184 => x"8cec0827",
          2185 => x"8b389816",
          2186 => x"08828cec",
          2187 => x"08268538",
          2188 => x"8258bd39",
          2189 => x"74733155",
          2190 => x"cb397352",
          2191 => x"7551f4d5",
          2192 => x"3f828cec",
          2193 => x"0898180c",
          2194 => x"7394180c",
          2195 => x"98170853",
          2196 => x"82587280",
          2197 => x"2e9a3885",
          2198 => x"39815894",
          2199 => x"3974892a",
          2200 => x"1398180c",
          2201 => x"7483ff06",
          2202 => x"16b4059c",
          2203 => x"180c8058",
          2204 => x"77828cec",
          2205 => x"0c8a3d0d",
          2206 => x"04f83d0d",
          2207 => x"7a700890",
          2208 => x"1208a005",
          2209 => x"595754f0",
          2210 => x"800a7727",
          2211 => x"8638800b",
          2212 => x"98150c98",
          2213 => x"14085384",
          2214 => x"5572802e",
          2215 => x"81cb3876",
          2216 => x"83ff0658",
          2217 => x"7781b538",
          2218 => x"81139815",
          2219 => x"0c941408",
          2220 => x"55749238",
          2221 => x"76852a88",
          2222 => x"17225653",
          2223 => x"74732681",
          2224 => x"9b3880c0",
          2225 => x"398a1622",
          2226 => x"ff057789",
          2227 => x"2a065372",
          2228 => x"818a3874",
          2229 => x"527351f3",
          2230 => x"e63f828c",
          2231 => x"ec085382",
          2232 => x"55810b82",
          2233 => x"8cec0827",
          2234 => x"80ff3881",
          2235 => x"55828cec",
          2236 => x"08ff2e80",
          2237 => x"f4389816",
          2238 => x"08828cec",
          2239 => x"082680ca",
          2240 => x"387b8a38",
          2241 => x"7798150c",
          2242 => x"845580dd",
          2243 => x"39941408",
          2244 => x"527351f9",
          2245 => x"863f828c",
          2246 => x"ec085387",
          2247 => x"55828cec",
          2248 => x"08802e80",
          2249 => x"c4388255",
          2250 => x"828cec08",
          2251 => x"812eba38",
          2252 => x"8155828c",
          2253 => x"ec08ff2e",
          2254 => x"b038828c",
          2255 => x"ec085275",
          2256 => x"51fbf33f",
          2257 => x"828cec08",
          2258 => x"a0387294",
          2259 => x"150c7252",
          2260 => x"7551f2c1",
          2261 => x"3f828cec",
          2262 => x"0898150c",
          2263 => x"7690150c",
          2264 => x"7716b405",
          2265 => x"9c150c80",
          2266 => x"5574828c",
          2267 => x"ec0c8a3d",
          2268 => x"0d04f73d",
          2269 => x"0d7b7d71",
          2270 => x"085b5b57",
          2271 => x"80527651",
          2272 => x"fcac3f82",
          2273 => x"8cec0854",
          2274 => x"828cec08",
          2275 => x"80ec3882",
          2276 => x"8cec0856",
          2277 => x"98170852",
          2278 => x"7851f083",
          2279 => x"3f828cec",
          2280 => x"0854828c",
          2281 => x"ec0880d2",
          2282 => x"38828cec",
          2283 => x"089c1808",
          2284 => x"70335154",
          2285 => x"587281e5",
          2286 => x"2e098106",
          2287 => x"83388158",
          2288 => x"828cec08",
          2289 => x"55728338",
          2290 => x"81557775",
          2291 => x"07537280",
          2292 => x"2e8e3881",
          2293 => x"1656757a",
          2294 => x"2e098106",
          2295 => x"8838a539",
          2296 => x"828cec08",
          2297 => x"56815276",
          2298 => x"51fd8e3f",
          2299 => x"828cec08",
          2300 => x"54828cec",
          2301 => x"08802eff",
          2302 => x"9b387384",
          2303 => x"2e098106",
          2304 => x"83388754",
          2305 => x"73828cec",
          2306 => x"0c8b3d0d",
          2307 => x"04fd3d0d",
          2308 => x"769a1152",
          2309 => x"54ebec3f",
          2310 => x"828cec08",
          2311 => x"83ffff06",
          2312 => x"76703351",
          2313 => x"53537183",
          2314 => x"2e098106",
          2315 => x"90389414",
          2316 => x"51ebd03f",
          2317 => x"828cec08",
          2318 => x"902b7307",
          2319 => x"5372828c",
          2320 => x"ec0c853d",
          2321 => x"0d04fc3d",
          2322 => x"0d777970",
          2323 => x"83ffff06",
          2324 => x"549a1253",
          2325 => x"5555ebed",
          2326 => x"3f767033",
          2327 => x"51537283",
          2328 => x"2e098106",
          2329 => x"8b387390",
          2330 => x"2a529415",
          2331 => x"51ebd63f",
          2332 => x"863d0d04",
          2333 => x"f73d0d7b",
          2334 => x"7d5b5584",
          2335 => x"75085a58",
          2336 => x"98150880",
          2337 => x"2e818a38",
          2338 => x"98150852",
          2339 => x"7851ee8f",
          2340 => x"3f828cec",
          2341 => x"0858828c",
          2342 => x"ec0880f5",
          2343 => x"389c1508",
          2344 => x"70335553",
          2345 => x"73863884",
          2346 => x"5880e639",
          2347 => x"8b133370",
          2348 => x"bf067081",
          2349 => x"ff065851",
          2350 => x"53728616",
          2351 => x"34828cec",
          2352 => x"08537381",
          2353 => x"e52e8338",
          2354 => x"815373ae",
          2355 => x"2ea93881",
          2356 => x"70740654",
          2357 => x"5772802e",
          2358 => x"9e38758f",
          2359 => x"2e993882",
          2360 => x"8cec0876",
          2361 => x"df065454",
          2362 => x"72882e09",
          2363 => x"81068338",
          2364 => x"7654737a",
          2365 => x"2ea03880",
          2366 => x"527451fa",
          2367 => x"fc3f828c",
          2368 => x"ec085882",
          2369 => x"8cec0889",
          2370 => x"38981508",
          2371 => x"fefa3886",
          2372 => x"39800b98",
          2373 => x"160c7782",
          2374 => x"8cec0c8b",
          2375 => x"3d0d04fb",
          2376 => x"3d0d7770",
          2377 => x"08575481",
          2378 => x"527351fc",
          2379 => x"c53f828c",
          2380 => x"ec085582",
          2381 => x"8cec08b4",
          2382 => x"38981408",
          2383 => x"527551ec",
          2384 => x"de3f828c",
          2385 => x"ec085582",
          2386 => x"8cec08a0",
          2387 => x"38a05382",
          2388 => x"8cec0852",
          2389 => x"9c140851",
          2390 => x"eadb3f8b",
          2391 => x"53a01452",
          2392 => x"9c140851",
          2393 => x"eaac3f81",
          2394 => x"0b831734",
          2395 => x"74828cec",
          2396 => x"0c873d0d",
          2397 => x"04fd3d0d",
          2398 => x"75700898",
          2399 => x"12085470",
          2400 => x"535553ec",
          2401 => x"9a3f828c",
          2402 => x"ec088d38",
          2403 => x"9c130853",
          2404 => x"e5733481",
          2405 => x"0b831534",
          2406 => x"853d0d04",
          2407 => x"fa3d0d78",
          2408 => x"7a575780",
          2409 => x"0b891734",
          2410 => x"98170880",
          2411 => x"2e818238",
          2412 => x"80708918",
          2413 => x"5555559c",
          2414 => x"17081470",
          2415 => x"33811656",
          2416 => x"515271a0",
          2417 => x"2ea83871",
          2418 => x"852e0981",
          2419 => x"06843881",
          2420 => x"e5527389",
          2421 => x"2e098106",
          2422 => x"8b38ae73",
          2423 => x"70810555",
          2424 => x"34811555",
          2425 => x"71737081",
          2426 => x"05553481",
          2427 => x"15558a74",
          2428 => x"27c53875",
          2429 => x"15880552",
          2430 => x"800b8113",
          2431 => x"349c1708",
          2432 => x"528b1233",
          2433 => x"8817349c",
          2434 => x"17089c11",
          2435 => x"5252e88a",
          2436 => x"3f828cec",
          2437 => x"08760c96",
          2438 => x"1251e7e7",
          2439 => x"3f828cec",
          2440 => x"08861723",
          2441 => x"981251e7",
          2442 => x"da3f828c",
          2443 => x"ec088417",
          2444 => x"23883d0d",
          2445 => x"04f33d0d",
          2446 => x"7f70085e",
          2447 => x"5b806170",
          2448 => x"33515555",
          2449 => x"73af2e83",
          2450 => x"38815573",
          2451 => x"80dc2e91",
          2452 => x"3874802e",
          2453 => x"8c38941d",
          2454 => x"08881c0c",
          2455 => x"aa398115",
          2456 => x"41806170",
          2457 => x"33565656",
          2458 => x"73af2e09",
          2459 => x"81068338",
          2460 => x"81567380",
          2461 => x"dc327030",
          2462 => x"70802578",
          2463 => x"07515154",
          2464 => x"73dc3873",
          2465 => x"881c0c60",
          2466 => x"70335154",
          2467 => x"739f2696",
          2468 => x"38ff800b",
          2469 => x"ab1c3480",
          2470 => x"527a51f6",
          2471 => x"913f828c",
          2472 => x"ec085585",
          2473 => x"9839913d",
          2474 => x"61a01d5c",
          2475 => x"5a5e8b53",
          2476 => x"a0527951",
          2477 => x"e7ff3f80",
          2478 => x"70595788",
          2479 => x"7933555c",
          2480 => x"73ae2e09",
          2481 => x"810680d4",
          2482 => x"38781870",
          2483 => x"33811a71",
          2484 => x"ae327030",
          2485 => x"709f2a73",
          2486 => x"82260751",
          2487 => x"51535a57",
          2488 => x"54738c38",
          2489 => x"79175475",
          2490 => x"74348117",
          2491 => x"57db3975",
          2492 => x"af327030",
          2493 => x"709f2a51",
          2494 => x"51547580",
          2495 => x"dc2e8c38",
          2496 => x"73802e87",
          2497 => x"3875a026",
          2498 => x"82bd3877",
          2499 => x"197e0ca4",
          2500 => x"54a07627",
          2501 => x"82bd38a0",
          2502 => x"5482b839",
          2503 => x"78187033",
          2504 => x"811a5a57",
          2505 => x"54a07627",
          2506 => x"81fc3875",
          2507 => x"af327030",
          2508 => x"7780dc32",
          2509 => x"70307280",
          2510 => x"25718025",
          2511 => x"07515156",
          2512 => x"51557380",
          2513 => x"2eac3884",
          2514 => x"39811858",
          2515 => x"80781a70",
          2516 => x"33515555",
          2517 => x"73af2e09",
          2518 => x"81068338",
          2519 => x"81557380",
          2520 => x"dc327030",
          2521 => x"70802577",
          2522 => x"07515154",
          2523 => x"73db3881",
          2524 => x"b53975ae",
          2525 => x"2e098106",
          2526 => x"83388154",
          2527 => x"767c2774",
          2528 => x"07547380",
          2529 => x"2ea2387b",
          2530 => x"8b327030",
          2531 => x"77ae3270",
          2532 => x"30728025",
          2533 => x"719f2a07",
          2534 => x"53515651",
          2535 => x"557481a7",
          2536 => x"3888578b",
          2537 => x"5cfef539",
          2538 => x"75982b54",
          2539 => x"7380258c",
          2540 => x"387580ff",
          2541 => x"0681fcbc",
          2542 => x"11335754",
          2543 => x"7551e6e1",
          2544 => x"3f828cec",
          2545 => x"08802eb2",
          2546 => x"38781870",
          2547 => x"33811a71",
          2548 => x"545a5654",
          2549 => x"e6d23f82",
          2550 => x"8cec0880",
          2551 => x"2e80e838",
          2552 => x"ff1c5476",
          2553 => x"742780df",
          2554 => x"38791754",
          2555 => x"75743481",
          2556 => x"177a1155",
          2557 => x"57747434",
          2558 => x"a7397552",
          2559 => x"81fbdc51",
          2560 => x"e5fe3f82",
          2561 => x"8cec08bf",
          2562 => x"38ff9f16",
          2563 => x"54739926",
          2564 => x"8938e016",
          2565 => x"7081ff06",
          2566 => x"57547917",
          2567 => x"54757434",
          2568 => x"811757fd",
          2569 => x"f7397719",
          2570 => x"7e0c7680",
          2571 => x"2e993879",
          2572 => x"33547381",
          2573 => x"e52e0981",
          2574 => x"06843885",
          2575 => x"7a348454",
          2576 => x"a076278f",
          2577 => x"388b3986",
          2578 => x"5581f239",
          2579 => x"845680f3",
          2580 => x"39805473",
          2581 => x"8b1b3480",
          2582 => x"7b085852",
          2583 => x"7a51f2ce",
          2584 => x"3f828cec",
          2585 => x"0856828c",
          2586 => x"ec0880d7",
          2587 => x"38981b08",
          2588 => x"527651e6",
          2589 => x"aa3f828c",
          2590 => x"ec085682",
          2591 => x"8cec0880",
          2592 => x"c2389c1b",
          2593 => x"08703355",
          2594 => x"5573802e",
          2595 => x"ffbe388b",
          2596 => x"1533bf06",
          2597 => x"5473861c",
          2598 => x"348b1533",
          2599 => x"70832a70",
          2600 => x"81065155",
          2601 => x"58739238",
          2602 => x"8b537952",
          2603 => x"7451e49f",
          2604 => x"3f828cec",
          2605 => x"08802e8b",
          2606 => x"3875527a",
          2607 => x"51f3ba3f",
          2608 => x"ff9f3975",
          2609 => x"ab1c3357",
          2610 => x"5574802e",
          2611 => x"bb387484",
          2612 => x"2e098106",
          2613 => x"80e73875",
          2614 => x"852a7081",
          2615 => x"0677822a",
          2616 => x"58515473",
          2617 => x"802e9638",
          2618 => x"75810654",
          2619 => x"73802efb",
          2620 => x"b538ff80",
          2621 => x"0bab1c34",
          2622 => x"805580c1",
          2623 => x"39758106",
          2624 => x"5473ba38",
          2625 => x"8555b639",
          2626 => x"75822a70",
          2627 => x"81065154",
          2628 => x"73ab3886",
          2629 => x"1b337084",
          2630 => x"2a708106",
          2631 => x"51555573",
          2632 => x"802ee138",
          2633 => x"901b0883",
          2634 => x"ff061db4",
          2635 => x"05527c51",
          2636 => x"f5db3f82",
          2637 => x"8cec0888",
          2638 => x"1c0cfaea",
          2639 => x"3974828c",
          2640 => x"ec0c8f3d",
          2641 => x"0d04f63d",
          2642 => x"0d7c5bff",
          2643 => x"7b087071",
          2644 => x"7355595c",
          2645 => x"55597380",
          2646 => x"2e81c638",
          2647 => x"75708105",
          2648 => x"573370a0",
          2649 => x"26525271",
          2650 => x"ba2e8d38",
          2651 => x"70ee3871",
          2652 => x"ba2e0981",
          2653 => x"0681a538",
          2654 => x"7333d011",
          2655 => x"7081ff06",
          2656 => x"51525370",
          2657 => x"89269138",
          2658 => x"82147381",
          2659 => x"ff06d005",
          2660 => x"56527176",
          2661 => x"2e80f738",
          2662 => x"800b81fc",
          2663 => x"ac595577",
          2664 => x"087a5557",
          2665 => x"76708105",
          2666 => x"58337470",
          2667 => x"81055633",
          2668 => x"ff9f1253",
          2669 => x"53537099",
          2670 => x"268938e0",
          2671 => x"137081ff",
          2672 => x"065451ff",
          2673 => x"9f125170",
          2674 => x"99268938",
          2675 => x"e0127081",
          2676 => x"ff065351",
          2677 => x"7230709f",
          2678 => x"2a515172",
          2679 => x"722e0981",
          2680 => x"06853870",
          2681 => x"ffbe3872",
          2682 => x"30747732",
          2683 => x"70307072",
          2684 => x"079f2a73",
          2685 => x"9f2a0753",
          2686 => x"54545170",
          2687 => x"802e8f38",
          2688 => x"81158419",
          2689 => x"59558375",
          2690 => x"25ff9438",
          2691 => x"8b397483",
          2692 => x"24863874",
          2693 => x"767c0c59",
          2694 => x"78518639",
          2695 => x"828d9c33",
          2696 => x"5170828c",
          2697 => x"ec0c8c3d",
          2698 => x"0d04fa3d",
          2699 => x"0d785680",
          2700 => x"0b831734",
          2701 => x"ff0bb017",
          2702 => x"0c795275",
          2703 => x"51e2e03f",
          2704 => x"8455828c",
          2705 => x"ec088180",
          2706 => x"3884b216",
          2707 => x"51dfb43f",
          2708 => x"828cec08",
          2709 => x"83ffff06",
          2710 => x"54835573",
          2711 => x"82d4d52e",
          2712 => x"09810680",
          2713 => x"e338800b",
          2714 => x"b4173356",
          2715 => x"577481e9",
          2716 => x"2e098106",
          2717 => x"83388157",
          2718 => x"7481eb32",
          2719 => x"70307080",
          2720 => x"25790751",
          2721 => x"5154738a",
          2722 => x"387481e8",
          2723 => x"2e098106",
          2724 => x"b5388353",
          2725 => x"81fbec52",
          2726 => x"80ea1651",
          2727 => x"e0b13f82",
          2728 => x"8cec0855",
          2729 => x"828cec08",
          2730 => x"802e9d38",
          2731 => x"855381fb",
          2732 => x"f0528186",
          2733 => x"1651e097",
          2734 => x"3f828cec",
          2735 => x"0855828c",
          2736 => x"ec08802e",
          2737 => x"83388255",
          2738 => x"74828cec",
          2739 => x"0c883d0d",
          2740 => x"04f23d0d",
          2741 => x"61028405",
          2742 => x"80cb0533",
          2743 => x"58558075",
          2744 => x"0c6051fc",
          2745 => x"e13f828c",
          2746 => x"ec08588b",
          2747 => x"56800b82",
          2748 => x"8cec0824",
          2749 => x"86fc3882",
          2750 => x"8cec0884",
          2751 => x"29828d88",
          2752 => x"05700855",
          2753 => x"538c5673",
          2754 => x"802e86e6",
          2755 => x"3873750c",
          2756 => x"7681fe06",
          2757 => x"74335457",
          2758 => x"72802eae",
          2759 => x"38811433",
          2760 => x"51d7ca3f",
          2761 => x"828cec08",
          2762 => x"81ff0670",
          2763 => x"81065455",
          2764 => x"72983876",
          2765 => x"802e86b8",
          2766 => x"3874822a",
          2767 => x"70810651",
          2768 => x"538a5672",
          2769 => x"86ac3886",
          2770 => x"a7398074",
          2771 => x"34778115",
          2772 => x"34815281",
          2773 => x"143351d7",
          2774 => x"b23f828c",
          2775 => x"ec0881ff",
          2776 => x"06708106",
          2777 => x"54558356",
          2778 => x"72868738",
          2779 => x"76802e8f",
          2780 => x"3874822a",
          2781 => x"70810651",
          2782 => x"538a5672",
          2783 => x"85f43880",
          2784 => x"70537452",
          2785 => x"5bfda33f",
          2786 => x"828cec08",
          2787 => x"81ff0657",
          2788 => x"76822e09",
          2789 => x"810680e2",
          2790 => x"388c3d74",
          2791 => x"56588356",
          2792 => x"83f61533",
          2793 => x"70585372",
          2794 => x"802e8d38",
          2795 => x"83fa1551",
          2796 => x"dce83f82",
          2797 => x"8cec0857",
          2798 => x"76787084",
          2799 => x"055a0cff",
          2800 => x"16901656",
          2801 => x"56758025",
          2802 => x"d738800b",
          2803 => x"8d3d5456",
          2804 => x"72708405",
          2805 => x"54085b83",
          2806 => x"577a802e",
          2807 => x"95387a52",
          2808 => x"7351fcc6",
          2809 => x"3f828cec",
          2810 => x"0881ff06",
          2811 => x"57817727",
          2812 => x"89388116",
          2813 => x"56837627",
          2814 => x"d7388156",
          2815 => x"76842e84",
          2816 => x"f1388d56",
          2817 => x"76812684",
          2818 => x"e938bf14",
          2819 => x"51dbf43f",
          2820 => x"828cec08",
          2821 => x"83ffff06",
          2822 => x"53728480",
          2823 => x"2e098106",
          2824 => x"84d03880",
          2825 => x"ca1451db",
          2826 => x"da3f828c",
          2827 => x"ec0883ff",
          2828 => x"ff065877",
          2829 => x"8d3880d8",
          2830 => x"1451dbde",
          2831 => x"3f828cec",
          2832 => x"0858779c",
          2833 => x"150c80c4",
          2834 => x"14338215",
          2835 => x"3480c414",
          2836 => x"33ff1170",
          2837 => x"81ff0651",
          2838 => x"54558d56",
          2839 => x"72812684",
          2840 => x"91387481",
          2841 => x"ff067871",
          2842 => x"2980c116",
          2843 => x"33525953",
          2844 => x"728a1523",
          2845 => x"72802e8b",
          2846 => x"38ff1373",
          2847 => x"06537280",
          2848 => x"2e86388d",
          2849 => x"5683eb39",
          2850 => x"80c51451",
          2851 => x"daf53f82",
          2852 => x"8cec0853",
          2853 => x"828cec08",
          2854 => x"88152372",
          2855 => x"8f06578d",
          2856 => x"567683ce",
          2857 => x"3880c714",
          2858 => x"51dad83f",
          2859 => x"828cec08",
          2860 => x"83ffff06",
          2861 => x"55748d38",
          2862 => x"80d41451",
          2863 => x"dadc3f82",
          2864 => x"8cec0855",
          2865 => x"80c21451",
          2866 => x"dab93f82",
          2867 => x"8cec0883",
          2868 => x"ffff0653",
          2869 => x"8d567280",
          2870 => x"2e839738",
          2871 => x"88142278",
          2872 => x"1471842a",
          2873 => x"055a5a78",
          2874 => x"75268386",
          2875 => x"388a1422",
          2876 => x"52747931",
          2877 => x"51ffb0be",
          2878 => x"3f828cec",
          2879 => x"0855828c",
          2880 => x"ec08802e",
          2881 => x"82ec3882",
          2882 => x"8cec0880",
          2883 => x"fffffff5",
          2884 => x"26833883",
          2885 => x"577483ff",
          2886 => x"f5268338",
          2887 => x"8257749f",
          2888 => x"f5268538",
          2889 => x"81578939",
          2890 => x"8d567680",
          2891 => x"2e82c338",
          2892 => x"82157098",
          2893 => x"160c7ba0",
          2894 => x"160c731c",
          2895 => x"70a4170c",
          2896 => x"7a1dac17",
          2897 => x"0c545576",
          2898 => x"832e0981",
          2899 => x"06af3880",
          2900 => x"de1451d9",
          2901 => x"ae3f828c",
          2902 => x"ec0883ff",
          2903 => x"ff06538d",
          2904 => x"5672828e",
          2905 => x"3879828a",
          2906 => x"3880e014",
          2907 => x"51d9ab3f",
          2908 => x"828cec08",
          2909 => x"a8150c74",
          2910 => x"822b53a2",
          2911 => x"398d5679",
          2912 => x"802e81ee",
          2913 => x"387713a8",
          2914 => x"150c7415",
          2915 => x"5376822e",
          2916 => x"8d387410",
          2917 => x"1570812a",
          2918 => x"76810605",
          2919 => x"515383ff",
          2920 => x"13892a53",
          2921 => x"8d56729c",
          2922 => x"15082681",
          2923 => x"c538ff0b",
          2924 => x"90150cff",
          2925 => x"0b8c150c",
          2926 => x"ff800b84",
          2927 => x"15347683",
          2928 => x"2e098106",
          2929 => x"81923880",
          2930 => x"e41451d8",
          2931 => x"b63f828c",
          2932 => x"ec0883ff",
          2933 => x"ff065372",
          2934 => x"812e0981",
          2935 => x"0680f938",
          2936 => x"811b5273",
          2937 => x"51dbb83f",
          2938 => x"828cec08",
          2939 => x"80ea3882",
          2940 => x"8cec0884",
          2941 => x"153484b2",
          2942 => x"1451d887",
          2943 => x"3f828cec",
          2944 => x"0883ffff",
          2945 => x"06537282",
          2946 => x"d4d52e09",
          2947 => x"810680c8",
          2948 => x"38b41451",
          2949 => x"d8843f82",
          2950 => x"8cec0884",
          2951 => x"8b85a4d2",
          2952 => x"2e098106",
          2953 => x"b3388498",
          2954 => x"1451d7ee",
          2955 => x"3f828cec",
          2956 => x"08868a85",
          2957 => x"e4f22e09",
          2958 => x"81069d38",
          2959 => x"849c1451",
          2960 => x"d7d83f82",
          2961 => x"8cec0890",
          2962 => x"150c84a0",
          2963 => x"1451d7ca",
          2964 => x"3f828cec",
          2965 => x"088c150c",
          2966 => x"76743482",
          2967 => x"8d982281",
          2968 => x"05537282",
          2969 => x"8d982372",
          2970 => x"86152380",
          2971 => x"0b94150c",
          2972 => x"80567582",
          2973 => x"8cec0c90",
          2974 => x"3d0d04fb",
          2975 => x"3d0d7754",
          2976 => x"89557380",
          2977 => x"2eb93873",
          2978 => x"08537280",
          2979 => x"2eb13872",
          2980 => x"33527180",
          2981 => x"2ea93886",
          2982 => x"13228415",
          2983 => x"22575271",
          2984 => x"762e0981",
          2985 => x"06993881",
          2986 => x"133351d0",
          2987 => x"c03f828c",
          2988 => x"ec088106",
          2989 => x"52718838",
          2990 => x"71740854",
          2991 => x"55833980",
          2992 => x"53787371",
          2993 => x"0c527482",
          2994 => x"8cec0c87",
          2995 => x"3d0d04fa",
          2996 => x"3d0d02ab",
          2997 => x"05337a58",
          2998 => x"893dfc05",
          2999 => x"5256f4e6",
          3000 => x"3f8b5480",
          3001 => x"0b828cec",
          3002 => x"0824bc38",
          3003 => x"828cec08",
          3004 => x"8429828d",
          3005 => x"88057008",
          3006 => x"55557380",
          3007 => x"2e843880",
          3008 => x"74347854",
          3009 => x"73802e84",
          3010 => x"38807434",
          3011 => x"78750c75",
          3012 => x"5475802e",
          3013 => x"92388053",
          3014 => x"893d7053",
          3015 => x"840551f7",
          3016 => x"b03f828c",
          3017 => x"ec085473",
          3018 => x"828cec0c",
          3019 => x"883d0d04",
          3020 => x"eb3d0d67",
          3021 => x"02840580",
          3022 => x"e7053359",
          3023 => x"59895478",
          3024 => x"802e84c8",
          3025 => x"3877bf06",
          3026 => x"7054983d",
          3027 => x"d0055399",
          3028 => x"3d840552",
          3029 => x"58f6fa3f",
          3030 => x"828cec08",
          3031 => x"55828cec",
          3032 => x"0884a438",
          3033 => x"7a5c6852",
          3034 => x"8c3d7052",
          3035 => x"56edc63f",
          3036 => x"828cec08",
          3037 => x"55828cec",
          3038 => x"08923802",
          3039 => x"80d70533",
          3040 => x"70982b55",
          3041 => x"57738025",
          3042 => x"83388655",
          3043 => x"779c0654",
          3044 => x"73802e81",
          3045 => x"ab387480",
          3046 => x"2e953874",
          3047 => x"842e0981",
          3048 => x"06aa3875",
          3049 => x"51eaf83f",
          3050 => x"828cec08",
          3051 => x"559e3902",
          3052 => x"b2053391",
          3053 => x"06547381",
          3054 => x"b8387782",
          3055 => x"2a708106",
          3056 => x"51547380",
          3057 => x"2e8e3888",
          3058 => x"5583bc39",
          3059 => x"77880758",
          3060 => x"7483b438",
          3061 => x"77832a70",
          3062 => x"81065154",
          3063 => x"73802e81",
          3064 => x"af386252",
          3065 => x"7a51e8a5",
          3066 => x"3f828cec",
          3067 => x"08568288",
          3068 => x"b20a5262",
          3069 => x"8e0551d4",
          3070 => x"ea3f6254",
          3071 => x"a00b8b15",
          3072 => x"34805362",
          3073 => x"527a51e8",
          3074 => x"bd3f8052",
          3075 => x"629c0551",
          3076 => x"d4d13f7a",
          3077 => x"54810b83",
          3078 => x"15347580",
          3079 => x"2e80f138",
          3080 => x"7ab01108",
          3081 => x"51548053",
          3082 => x"7552973d",
          3083 => x"d40551dd",
          3084 => x"be3f828c",
          3085 => x"ec085582",
          3086 => x"8cec0882",
          3087 => x"ca38b739",
          3088 => x"7482c438",
          3089 => x"02b20533",
          3090 => x"70842a70",
          3091 => x"81065155",
          3092 => x"5673802e",
          3093 => x"86388455",
          3094 => x"82ad3977",
          3095 => x"812a7081",
          3096 => x"06515473",
          3097 => x"802ea938",
          3098 => x"75810654",
          3099 => x"73802ea0",
          3100 => x"38875582",
          3101 => x"92397352",
          3102 => x"7a51d6a3",
          3103 => x"3f828cec",
          3104 => x"087bff18",
          3105 => x"8c120c55",
          3106 => x"55828cec",
          3107 => x"0881f838",
          3108 => x"77832a70",
          3109 => x"81065154",
          3110 => x"73802e86",
          3111 => x"387780c0",
          3112 => x"07587ab0",
          3113 => x"1108a01b",
          3114 => x"0c63a41b",
          3115 => x"0c635370",
          3116 => x"5257e6d9",
          3117 => x"3f828cec",
          3118 => x"08828cec",
          3119 => x"08881b0c",
          3120 => x"639c0552",
          3121 => x"5ad2d33f",
          3122 => x"828cec08",
          3123 => x"828cec08",
          3124 => x"8c1b0c77",
          3125 => x"7a0c5686",
          3126 => x"1722841a",
          3127 => x"2377901a",
          3128 => x"34800b91",
          3129 => x"1a34800b",
          3130 => x"9c1a0c80",
          3131 => x"0b941a0c",
          3132 => x"77852a70",
          3133 => x"81065154",
          3134 => x"73802e81",
          3135 => x"8d38828c",
          3136 => x"ec08802e",
          3137 => x"81843882",
          3138 => x"8cec0894",
          3139 => x"1a0c8a17",
          3140 => x"2270892b",
          3141 => x"7b525957",
          3142 => x"a8397652",
          3143 => x"7851d79f",
          3144 => x"3f828cec",
          3145 => x"0857828c",
          3146 => x"ec088126",
          3147 => x"83388255",
          3148 => x"828cec08",
          3149 => x"ff2e0981",
          3150 => x"06833879",
          3151 => x"55757831",
          3152 => x"56743070",
          3153 => x"76078025",
          3154 => x"51547776",
          3155 => x"278a3881",
          3156 => x"70750655",
          3157 => x"5a73c338",
          3158 => x"76981a0c",
          3159 => x"74a93875",
          3160 => x"83ff0654",
          3161 => x"73802ea2",
          3162 => x"3876527a",
          3163 => x"51d6a63f",
          3164 => x"828cec08",
          3165 => x"85388255",
          3166 => x"8e397589",
          3167 => x"2a828cec",
          3168 => x"08059c1a",
          3169 => x"0c843980",
          3170 => x"790c7454",
          3171 => x"73828cec",
          3172 => x"0c973d0d",
          3173 => x"04f23d0d",
          3174 => x"60636564",
          3175 => x"40405d59",
          3176 => x"807e0c90",
          3177 => x"3dfc0552",
          3178 => x"7851f9cf",
          3179 => x"3f828cec",
          3180 => x"0855828c",
          3181 => x"ec088a38",
          3182 => x"91193355",
          3183 => x"74802e86",
          3184 => x"38745682",
          3185 => x"c4399019",
          3186 => x"33810655",
          3187 => x"87567480",
          3188 => x"2e82b638",
          3189 => x"9539820b",
          3190 => x"911a3482",
          3191 => x"5682aa39",
          3192 => x"810b911a",
          3193 => x"34815682",
          3194 => x"a0398c19",
          3195 => x"08941a08",
          3196 => x"3155747c",
          3197 => x"27833874",
          3198 => x"5c7b802e",
          3199 => x"82893894",
          3200 => x"19087083",
          3201 => x"ff065656",
          3202 => x"7481b238",
          3203 => x"7e8a1122",
          3204 => x"ff057789",
          3205 => x"2a065b55",
          3206 => x"79a83875",
          3207 => x"87388819",
          3208 => x"08558f39",
          3209 => x"98190852",
          3210 => x"7851d593",
          3211 => x"3f828cec",
          3212 => x"08558175",
          3213 => x"27ff9f38",
          3214 => x"74ff2eff",
          3215 => x"a3387498",
          3216 => x"1a0c9819",
          3217 => x"08527e51",
          3218 => x"d4cb3f82",
          3219 => x"8cec0880",
          3220 => x"2eff8338",
          3221 => x"828cec08",
          3222 => x"1a7c892a",
          3223 => x"59577780",
          3224 => x"2e80d638",
          3225 => x"771a7f8a",
          3226 => x"1122585c",
          3227 => x"55757527",
          3228 => x"8538757a",
          3229 => x"31587754",
          3230 => x"76537c52",
          3231 => x"811b3351",
          3232 => x"ca883f82",
          3233 => x"8cec08fe",
          3234 => x"d7387e83",
          3235 => x"11335656",
          3236 => x"74802e9f",
          3237 => x"38b01608",
          3238 => x"77315574",
          3239 => x"78279438",
          3240 => x"848053b4",
          3241 => x"1652b016",
          3242 => x"08773189",
          3243 => x"2b7d0551",
          3244 => x"cfe03f77",
          3245 => x"892b56b9",
          3246 => x"39769c1a",
          3247 => x"0c941908",
          3248 => x"83ff0684",
          3249 => x"80713157",
          3250 => x"557b7627",
          3251 => x"83387b56",
          3252 => x"9c190852",
          3253 => x"7e51d1c7",
          3254 => x"3f828cec",
          3255 => x"08fe8138",
          3256 => x"75539419",
          3257 => x"0883ff06",
          3258 => x"1fb40552",
          3259 => x"7c51cfa2",
          3260 => x"3f7b7631",
          3261 => x"7e08177f",
          3262 => x"0c761e94",
          3263 => x"1b081894",
          3264 => x"1c0c5e5c",
          3265 => x"fdf33980",
          3266 => x"5675828c",
          3267 => x"ec0c903d",
          3268 => x"0d04f23d",
          3269 => x"0d606365",
          3270 => x"6440405d",
          3271 => x"58807e0c",
          3272 => x"903dfc05",
          3273 => x"527751f6",
          3274 => x"d23f828c",
          3275 => x"ec085582",
          3276 => x"8cec088a",
          3277 => x"38911833",
          3278 => x"5574802e",
          3279 => x"86387456",
          3280 => x"83b83990",
          3281 => x"18337081",
          3282 => x"2a708106",
          3283 => x"51565687",
          3284 => x"5674802e",
          3285 => x"83a43895",
          3286 => x"39820b91",
          3287 => x"19348256",
          3288 => x"83983981",
          3289 => x"0b911934",
          3290 => x"8156838e",
          3291 => x"39941808",
          3292 => x"7c115656",
          3293 => x"74762784",
          3294 => x"3875095c",
          3295 => x"7b802e82",
          3296 => x"ec389418",
          3297 => x"087083ff",
          3298 => x"06565674",
          3299 => x"81fd387e",
          3300 => x"8a1122ff",
          3301 => x"0577892a",
          3302 => x"065c557a",
          3303 => x"bf38758c",
          3304 => x"38881808",
          3305 => x"55749c38",
          3306 => x"7a528539",
          3307 => x"98180852",
          3308 => x"7751d7e7",
          3309 => x"3f828cec",
          3310 => x"0855828c",
          3311 => x"ec08802e",
          3312 => x"82ab3874",
          3313 => x"812eff91",
          3314 => x"3874ff2e",
          3315 => x"ff953874",
          3316 => x"98190c88",
          3317 => x"18088538",
          3318 => x"7488190c",
          3319 => x"7e55b015",
          3320 => x"089c1908",
          3321 => x"2e098106",
          3322 => x"8d387451",
          3323 => x"cec13f82",
          3324 => x"8cec08fe",
          3325 => x"ee389818",
          3326 => x"08527e51",
          3327 => x"d1973f82",
          3328 => x"8cec0880",
          3329 => x"2efed238",
          3330 => x"828cec08",
          3331 => x"1b7c892a",
          3332 => x"5a577880",
          3333 => x"2e80d538",
          3334 => x"781b7f8a",
          3335 => x"1122585b",
          3336 => x"55757527",
          3337 => x"8538757b",
          3338 => x"31597854",
          3339 => x"76537c52",
          3340 => x"811a3351",
          3341 => x"c8be3f82",
          3342 => x"8cec08fe",
          3343 => x"a6387eb0",
          3344 => x"11087831",
          3345 => x"56567479",
          3346 => x"279b3884",
          3347 => x"8053b016",
          3348 => x"08773189",
          3349 => x"2b7d0552",
          3350 => x"b41651cc",
          3351 => x"b53f7e55",
          3352 => x"800b8316",
          3353 => x"3478892b",
          3354 => x"5680db39",
          3355 => x"8c180894",
          3356 => x"19082693",
          3357 => x"387e51cd",
          3358 => x"b63f828c",
          3359 => x"ec08fde3",
          3360 => x"387e77b0",
          3361 => x"120c5576",
          3362 => x"9c190c94",
          3363 => x"180883ff",
          3364 => x"06848071",
          3365 => x"3157557b",
          3366 => x"76278338",
          3367 => x"7b569c18",
          3368 => x"08527e51",
          3369 => x"cdf93f82",
          3370 => x"8cec08fd",
          3371 => x"b6387553",
          3372 => x"7c529418",
          3373 => x"0883ff06",
          3374 => x"1fb40551",
          3375 => x"cbd43f7e",
          3376 => x"55810b83",
          3377 => x"16347b76",
          3378 => x"317e0817",
          3379 => x"7f0c761e",
          3380 => x"941a0818",
          3381 => x"70941c0c",
          3382 => x"8c1b0858",
          3383 => x"585e5c74",
          3384 => x"76278338",
          3385 => x"7555748c",
          3386 => x"190cfd90",
          3387 => x"39901833",
          3388 => x"80c00755",
          3389 => x"74901934",
          3390 => x"80567582",
          3391 => x"8cec0c90",
          3392 => x"3d0d04f8",
          3393 => x"3d0d7a8b",
          3394 => x"3dfc0553",
          3395 => x"705256f2",
          3396 => x"ea3f828c",
          3397 => x"ec085782",
          3398 => x"8cec0880",
          3399 => x"fb389016",
          3400 => x"3370862a",
          3401 => x"70810651",
          3402 => x"55557380",
          3403 => x"2e80e938",
          3404 => x"a0160852",
          3405 => x"7851cce7",
          3406 => x"3f828cec",
          3407 => x"0857828c",
          3408 => x"ec0880d4",
          3409 => x"38a41608",
          3410 => x"8b1133a0",
          3411 => x"07555573",
          3412 => x"8b163488",
          3413 => x"16085374",
          3414 => x"52750851",
          3415 => x"dde83f8c",
          3416 => x"1608529c",
          3417 => x"1551c9fb",
          3418 => x"3f8288b2",
          3419 => x"0a529615",
          3420 => x"51c9f03f",
          3421 => x"76529215",
          3422 => x"51c9ca3f",
          3423 => x"7854810b",
          3424 => x"83153478",
          3425 => x"51ccdf3f",
          3426 => x"828cec08",
          3427 => x"90173381",
          3428 => x"bf065557",
          3429 => x"73901734",
          3430 => x"76828cec",
          3431 => x"0c8a3d0d",
          3432 => x"04fc3d0d",
          3433 => x"76705254",
          3434 => x"fed93f82",
          3435 => x"8cec0853",
          3436 => x"828cec08",
          3437 => x"9c38863d",
          3438 => x"fc055273",
          3439 => x"51f1bc3f",
          3440 => x"828cec08",
          3441 => x"53828cec",
          3442 => x"08873882",
          3443 => x"8cec0874",
          3444 => x"0c72828c",
          3445 => x"ec0c863d",
          3446 => x"0d04ff3d",
          3447 => x"0d843d51",
          3448 => x"e6e43f8b",
          3449 => x"52800b82",
          3450 => x"8cec0824",
          3451 => x"8b38828c",
          3452 => x"ec08828d",
          3453 => x"9c348052",
          3454 => x"71828cec",
          3455 => x"0c833d0d",
          3456 => x"04ef3d0d",
          3457 => x"8053933d",
          3458 => x"d0055294",
          3459 => x"3d51e9c1",
          3460 => x"3f828cec",
          3461 => x"0855828c",
          3462 => x"ec0880e0",
          3463 => x"38765863",
          3464 => x"52933dd4",
          3465 => x"0551e08d",
          3466 => x"3f828cec",
          3467 => x"0855828c",
          3468 => x"ec08bc38",
          3469 => x"0280c705",
          3470 => x"3370982b",
          3471 => x"55567380",
          3472 => x"25893876",
          3473 => x"7a94120c",
          3474 => x"54b23902",
          3475 => x"a2053370",
          3476 => x"842a7081",
          3477 => x"06515556",
          3478 => x"73802e9e",
          3479 => x"38767f53",
          3480 => x"705254db",
          3481 => x"a83f828c",
          3482 => x"ec089415",
          3483 => x"0c8e3982",
          3484 => x"8cec0884",
          3485 => x"2e098106",
          3486 => x"83388555",
          3487 => x"74828cec",
          3488 => x"0c933d0d",
          3489 => x"04e43d0d",
          3490 => x"6f6f5b5b",
          3491 => x"807a3480",
          3492 => x"539e3dff",
          3493 => x"b805529f",
          3494 => x"3d51e8b5",
          3495 => x"3f828cec",
          3496 => x"0857828c",
          3497 => x"ec0882fc",
          3498 => x"387b437a",
          3499 => x"7c941108",
          3500 => x"47555864",
          3501 => x"5473802e",
          3502 => x"81ed38a0",
          3503 => x"52933d70",
          3504 => x"5255d5ea",
          3505 => x"3f828cec",
          3506 => x"0857828c",
          3507 => x"ec0882d4",
          3508 => x"3868527b",
          3509 => x"51c9c83f",
          3510 => x"828cec08",
          3511 => x"57828cec",
          3512 => x"0882c138",
          3513 => x"69527b51",
          3514 => x"daa33f82",
          3515 => x"8cec0845",
          3516 => x"76527451",
          3517 => x"d5b83f82",
          3518 => x"8cec0857",
          3519 => x"828cec08",
          3520 => x"82a23880",
          3521 => x"527451da",
          3522 => x"eb3f828c",
          3523 => x"ec085782",
          3524 => x"8cec08a4",
          3525 => x"3869527b",
          3526 => x"51d9f23f",
          3527 => x"73828cec",
          3528 => x"082ea638",
          3529 => x"76527451",
          3530 => x"d6cf3f82",
          3531 => x"8cec0857",
          3532 => x"828cec08",
          3533 => x"802ecc38",
          3534 => x"76842e09",
          3535 => x"81068638",
          3536 => x"825781e0",
          3537 => x"397681dc",
          3538 => x"389e3dff",
          3539 => x"bc055274",
          3540 => x"51dcc93f",
          3541 => x"76903d78",
          3542 => x"11811133",
          3543 => x"51565a56",
          3544 => x"73802e91",
          3545 => x"3802b905",
          3546 => x"55811681",
          3547 => x"16703356",
          3548 => x"565673f5",
          3549 => x"38811654",
          3550 => x"73782681",
          3551 => x"90387580",
          3552 => x"2e993878",
          3553 => x"16810555",
          3554 => x"ff186f11",
          3555 => x"ff18ff18",
          3556 => x"58585558",
          3557 => x"74337434",
          3558 => x"75ee38ff",
          3559 => x"186f1155",
          3560 => x"58af7434",
          3561 => x"fe8d3977",
          3562 => x"7b2e0981",
          3563 => x"068a38ff",
          3564 => x"186f1155",
          3565 => x"58af7434",
          3566 => x"800b828d",
          3567 => x"9c337084",
          3568 => x"2981fcac",
          3569 => x"05700870",
          3570 => x"33525c56",
          3571 => x"56567376",
          3572 => x"2e8d3881",
          3573 => x"16701a70",
          3574 => x"33515556",
          3575 => x"73f53882",
          3576 => x"16547378",
          3577 => x"26a73880",
          3578 => x"55747627",
          3579 => x"91387419",
          3580 => x"5473337a",
          3581 => x"7081055c",
          3582 => x"34811555",
          3583 => x"ec39ba7a",
          3584 => x"7081055c",
          3585 => x"3474ff2e",
          3586 => x"09810685",
          3587 => x"38915794",
          3588 => x"396e1881",
          3589 => x"19595473",
          3590 => x"337a7081",
          3591 => x"055c347a",
          3592 => x"7826ee38",
          3593 => x"807a3476",
          3594 => x"828cec0c",
          3595 => x"9e3d0d04",
          3596 => x"f73d0d7b",
          3597 => x"7d8d3dfc",
          3598 => x"05547153",
          3599 => x"5755ecbb",
          3600 => x"3f828cec",
          3601 => x"0853828c",
          3602 => x"ec0882fa",
          3603 => x"38911533",
          3604 => x"537282f2",
          3605 => x"388c1508",
          3606 => x"54737627",
          3607 => x"92389015",
          3608 => x"3370812a",
          3609 => x"70810651",
          3610 => x"54577283",
          3611 => x"38735694",
          3612 => x"15085480",
          3613 => x"7094170c",
          3614 => x"5875782e",
          3615 => x"82973879",
          3616 => x"8a112270",
          3617 => x"892b5951",
          3618 => x"5373782e",
          3619 => x"b7387652",
          3620 => x"ff1651ff",
          3621 => x"99a03f82",
          3622 => x"8cec08ff",
          3623 => x"15785470",
          3624 => x"535553ff",
          3625 => x"99903f82",
          3626 => x"8cec0873",
          3627 => x"26963876",
          3628 => x"30707506",
          3629 => x"7094180c",
          3630 => x"77713198",
          3631 => x"18085758",
          3632 => x"5153b139",
          3633 => x"88150854",
          3634 => x"73a63873",
          3635 => x"527451cd",
          3636 => x"ca3f828c",
          3637 => x"ec085482",
          3638 => x"8cec0881",
          3639 => x"2e819a38",
          3640 => x"828cec08",
          3641 => x"ff2e819b",
          3642 => x"38828cec",
          3643 => x"0888160c",
          3644 => x"7398160c",
          3645 => x"73802e81",
          3646 => x"9c387676",
          3647 => x"2780dc38",
          3648 => x"75773194",
          3649 => x"16081894",
          3650 => x"170c9016",
          3651 => x"3370812a",
          3652 => x"70810651",
          3653 => x"555a5672",
          3654 => x"802e9a38",
          3655 => x"73527451",
          3656 => x"ccf93f82",
          3657 => x"8cec0854",
          3658 => x"828cec08",
          3659 => x"9438828c",
          3660 => x"ec0856a7",
          3661 => x"39735274",
          3662 => x"51c7843f",
          3663 => x"828cec08",
          3664 => x"5473ff2e",
          3665 => x"be388174",
          3666 => x"27af3879",
          3667 => x"53739814",
          3668 => x"0827a638",
          3669 => x"7398160c",
          3670 => x"ffa03994",
          3671 => x"15081694",
          3672 => x"160c7583",
          3673 => x"ff065372",
          3674 => x"802eaa38",
          3675 => x"73527951",
          3676 => x"c6a33f82",
          3677 => x"8cec0894",
          3678 => x"38820b91",
          3679 => x"16348253",
          3680 => x"80c43981",
          3681 => x"0b911634",
          3682 => x"8153bb39",
          3683 => x"75892a82",
          3684 => x"8cec0805",
          3685 => x"58941508",
          3686 => x"548c1508",
          3687 => x"74279038",
          3688 => x"738c160c",
          3689 => x"90153380",
          3690 => x"c0075372",
          3691 => x"90163473",
          3692 => x"83ff0653",
          3693 => x"72802e8c",
          3694 => x"38779c16",
          3695 => x"082e8538",
          3696 => x"779c160c",
          3697 => x"80537282",
          3698 => x"8cec0c8b",
          3699 => x"3d0d04f9",
          3700 => x"3d0d7956",
          3701 => x"89547580",
          3702 => x"2e818a38",
          3703 => x"8053893d",
          3704 => x"fc05528a",
          3705 => x"3d840551",
          3706 => x"e1e73f82",
          3707 => x"8cec0855",
          3708 => x"828cec08",
          3709 => x"80ea3877",
          3710 => x"760c7a52",
          3711 => x"7551d8b5",
          3712 => x"3f828cec",
          3713 => x"0855828c",
          3714 => x"ec0880c3",
          3715 => x"38ab1633",
          3716 => x"70982b55",
          3717 => x"57807424",
          3718 => x"a2388616",
          3719 => x"3370842a",
          3720 => x"70810651",
          3721 => x"55577380",
          3722 => x"2ead389c",
          3723 => x"16085277",
          3724 => x"51d3da3f",
          3725 => x"828cec08",
          3726 => x"88170c77",
          3727 => x"54861422",
          3728 => x"84172374",
          3729 => x"527551ce",
          3730 => x"e53f828c",
          3731 => x"ec085574",
          3732 => x"842e0981",
          3733 => x"06853885",
          3734 => x"55863974",
          3735 => x"802e8438",
          3736 => x"80760c74",
          3737 => x"5473828c",
          3738 => x"ec0c893d",
          3739 => x"0d04fc3d",
          3740 => x"0d76873d",
          3741 => x"fc055370",
          3742 => x"5253e7ff",
          3743 => x"3f828cec",
          3744 => x"08873882",
          3745 => x"8cec0873",
          3746 => x"0c863d0d",
          3747 => x"04fb3d0d",
          3748 => x"7779893d",
          3749 => x"fc055471",
          3750 => x"535654e7",
          3751 => x"de3f828c",
          3752 => x"ec085382",
          3753 => x"8cec0880",
          3754 => x"df387493",
          3755 => x"38828cec",
          3756 => x"08527351",
          3757 => x"cdf83f82",
          3758 => x"8cec0853",
          3759 => x"80ca3982",
          3760 => x"8cec0852",
          3761 => x"7351d3ac",
          3762 => x"3f828cec",
          3763 => x"0853828c",
          3764 => x"ec08842e",
          3765 => x"09810685",
          3766 => x"38805387",
          3767 => x"39828cec",
          3768 => x"08a63874",
          3769 => x"527351d5",
          3770 => x"b33f7252",
          3771 => x"7351cf89",
          3772 => x"3f828cec",
          3773 => x"08843270",
          3774 => x"30707207",
          3775 => x"9f2c7082",
          3776 => x"8cec0806",
          3777 => x"51515454",
          3778 => x"72828cec",
          3779 => x"0c873d0d",
          3780 => x"04ee3d0d",
          3781 => x"65578053",
          3782 => x"893d7053",
          3783 => x"963d5256",
          3784 => x"dfaf3f82",
          3785 => x"8cec0855",
          3786 => x"828cec08",
          3787 => x"b2386452",
          3788 => x"7551d681",
          3789 => x"3f828cec",
          3790 => x"0855828c",
          3791 => x"ec08a038",
          3792 => x"0280cb05",
          3793 => x"3370982b",
          3794 => x"55587380",
          3795 => x"25853886",
          3796 => x"558d3976",
          3797 => x"802e8838",
          3798 => x"76527551",
          3799 => x"d4be3f74",
          3800 => x"828cec0c",
          3801 => x"943d0d04",
          3802 => x"f03d0d63",
          3803 => x"65555c80",
          3804 => x"53923dec",
          3805 => x"0552933d",
          3806 => x"51ded63f",
          3807 => x"828cec08",
          3808 => x"5b828cec",
          3809 => x"08828038",
          3810 => x"7c740c73",
          3811 => x"08981108",
          3812 => x"fe119013",
          3813 => x"08595658",
          3814 => x"55757426",
          3815 => x"9138757c",
          3816 => x"0c81e439",
          3817 => x"815b81cc",
          3818 => x"39825b81",
          3819 => x"c739828c",
          3820 => x"ec087533",
          3821 => x"55597381",
          3822 => x"2e098106",
          3823 => x"bf388275",
          3824 => x"5f577652",
          3825 => x"923df005",
          3826 => x"51c1f43f",
          3827 => x"828cec08",
          3828 => x"ff2ed138",
          3829 => x"828cec08",
          3830 => x"812ece38",
          3831 => x"828cec08",
          3832 => x"3070828c",
          3833 => x"ec080780",
          3834 => x"257a0581",
          3835 => x"197f5359",
          3836 => x"5a549814",
          3837 => x"087726ca",
          3838 => x"3880f939",
          3839 => x"a4150882",
          3840 => x"8cec0857",
          3841 => x"58759838",
          3842 => x"77528118",
          3843 => x"7d5258ff",
          3844 => x"bf8d3f82",
          3845 => x"8cec085b",
          3846 => x"828cec08",
          3847 => x"80d6387c",
          3848 => x"70337712",
          3849 => x"ff1a5d52",
          3850 => x"56547482",
          3851 => x"2e098106",
          3852 => x"9e38b414",
          3853 => x"51ffbbcb",
          3854 => x"3f828cec",
          3855 => x"0883ffff",
          3856 => x"06703070",
          3857 => x"80251b82",
          3858 => x"19595b51",
          3859 => x"549b39b4",
          3860 => x"1451ffbb",
          3861 => x"c53f828c",
          3862 => x"ec08f00a",
          3863 => x"06703070",
          3864 => x"80251b84",
          3865 => x"19595b51",
          3866 => x"547583ff",
          3867 => x"067a5856",
          3868 => x"79ff9238",
          3869 => x"787c0c7c",
          3870 => x"7990120c",
          3871 => x"84113381",
          3872 => x"07565474",
          3873 => x"8415347a",
          3874 => x"828cec0c",
          3875 => x"923d0d04",
          3876 => x"f93d0d79",
          3877 => x"8a3dfc05",
          3878 => x"53705257",
          3879 => x"e3dd3f82",
          3880 => x"8cec0856",
          3881 => x"828cec08",
          3882 => x"81a83891",
          3883 => x"17335675",
          3884 => x"81a03890",
          3885 => x"17337081",
          3886 => x"2a708106",
          3887 => x"51555587",
          3888 => x"5573802e",
          3889 => x"818e3894",
          3890 => x"17085473",
          3891 => x"8c180827",
          3892 => x"81803873",
          3893 => x"9b38828c",
          3894 => x"ec085388",
          3895 => x"17085276",
          3896 => x"51c48c3f",
          3897 => x"828cec08",
          3898 => x"7488190c",
          3899 => x"5680c939",
          3900 => x"98170852",
          3901 => x"7651ffbf",
          3902 => x"c63f828c",
          3903 => x"ec08ff2e",
          3904 => x"09810683",
          3905 => x"38815682",
          3906 => x"8cec0881",
          3907 => x"2e098106",
          3908 => x"85388256",
          3909 => x"a33975a0",
          3910 => x"38775482",
          3911 => x"8cec0898",
          3912 => x"15082794",
          3913 => x"38981708",
          3914 => x"53828cec",
          3915 => x"08527651",
          3916 => x"c3bd3f82",
          3917 => x"8cec0856",
          3918 => x"9417088c",
          3919 => x"180c9017",
          3920 => x"3380c007",
          3921 => x"54739018",
          3922 => x"3475802e",
          3923 => x"85387591",
          3924 => x"18347555",
          3925 => x"74828cec",
          3926 => x"0c893d0d",
          3927 => x"04e23d0d",
          3928 => x"8253a03d",
          3929 => x"ffa40552",
          3930 => x"a13d51da",
          3931 => x"e43f828c",
          3932 => x"ec085582",
          3933 => x"8cec0881",
          3934 => x"f5387845",
          3935 => x"a13d0852",
          3936 => x"953d7052",
          3937 => x"58d1ae3f",
          3938 => x"828cec08",
          3939 => x"55828cec",
          3940 => x"0881db38",
          3941 => x"0280fb05",
          3942 => x"3370852a",
          3943 => x"70810651",
          3944 => x"55568655",
          3945 => x"7381c738",
          3946 => x"75982b54",
          3947 => x"80742481",
          3948 => x"bd380280",
          3949 => x"d6053370",
          3950 => x"81065854",
          3951 => x"87557681",
          3952 => x"ad386b52",
          3953 => x"7851ccc5",
          3954 => x"3f828cec",
          3955 => x"0874842a",
          3956 => x"70810651",
          3957 => x"55567380",
          3958 => x"2e80d438",
          3959 => x"7854828c",
          3960 => x"ec089415",
          3961 => x"082e8186",
          3962 => x"38735a82",
          3963 => x"8cec085c",
          3964 => x"76528a3d",
          3965 => x"705254c7",
          3966 => x"b53f828c",
          3967 => x"ec085582",
          3968 => x"8cec0880",
          3969 => x"e938828c",
          3970 => x"ec085273",
          3971 => x"51cce53f",
          3972 => x"828cec08",
          3973 => x"55828cec",
          3974 => x"08863887",
          3975 => x"5580cf39",
          3976 => x"828cec08",
          3977 => x"842e8838",
          3978 => x"828cec08",
          3979 => x"80c03877",
          3980 => x"51cec23f",
          3981 => x"828cec08",
          3982 => x"828cec08",
          3983 => x"3070828c",
          3984 => x"ec080780",
          3985 => x"25515555",
          3986 => x"75802e94",
          3987 => x"3873802e",
          3988 => x"8f388053",
          3989 => x"75527751",
          3990 => x"c1953f82",
          3991 => x"8cec0855",
          3992 => x"748c3878",
          3993 => x"51ffbafe",
          3994 => x"3f828cec",
          3995 => x"08557482",
          3996 => x"8cec0ca0",
          3997 => x"3d0d04e9",
          3998 => x"3d0d8253",
          3999 => x"993dc005",
          4000 => x"529a3d51",
          4001 => x"d8cb3f82",
          4002 => x"8cec0854",
          4003 => x"828cec08",
          4004 => x"82b03878",
          4005 => x"5e69528e",
          4006 => x"3d705258",
          4007 => x"cf973f82",
          4008 => x"8cec0854",
          4009 => x"828cec08",
          4010 => x"86388854",
          4011 => x"82943982",
          4012 => x"8cec0884",
          4013 => x"2e098106",
          4014 => x"82883802",
          4015 => x"80df0533",
          4016 => x"70852a81",
          4017 => x"06515586",
          4018 => x"547481f6",
          4019 => x"38785a74",
          4020 => x"528a3d70",
          4021 => x"5257c1c3",
          4022 => x"3f828cec",
          4023 => x"08755556",
          4024 => x"828cec08",
          4025 => x"83388754",
          4026 => x"828cec08",
          4027 => x"812e0981",
          4028 => x"06833882",
          4029 => x"54828cec",
          4030 => x"08ff2e09",
          4031 => x"81068638",
          4032 => x"815481b4",
          4033 => x"397381b0",
          4034 => x"38828cec",
          4035 => x"08527851",
          4036 => x"c4a43f82",
          4037 => x"8cec0854",
          4038 => x"828cec08",
          4039 => x"819a388b",
          4040 => x"53a052b4",
          4041 => x"1951ffb7",
          4042 => x"8c3f7854",
          4043 => x"ae0bb415",
          4044 => x"34785490",
          4045 => x"0bbf1534",
          4046 => x"8288b20a",
          4047 => x"5280ca19",
          4048 => x"51ffb69f",
          4049 => x"3f755378",
          4050 => x"b4115351",
          4051 => x"c9f83fa0",
          4052 => x"5378b411",
          4053 => x"5380d405",
          4054 => x"51ffb6b6",
          4055 => x"3f7854ae",
          4056 => x"0b80d515",
          4057 => x"347f5378",
          4058 => x"80d41153",
          4059 => x"51c9d73f",
          4060 => x"7854810b",
          4061 => x"83153477",
          4062 => x"51cba43f",
          4063 => x"828cec08",
          4064 => x"54828cec",
          4065 => x"08b23882",
          4066 => x"88b20a52",
          4067 => x"64960551",
          4068 => x"ffb5d03f",
          4069 => x"75536452",
          4070 => x"7851c9aa",
          4071 => x"3f645490",
          4072 => x"0b8b1534",
          4073 => x"7854810b",
          4074 => x"83153478",
          4075 => x"51ffb8b6",
          4076 => x"3f828cec",
          4077 => x"08548b39",
          4078 => x"80537552",
          4079 => x"7651ffbe",
          4080 => x"ae3f7382",
          4081 => x"8cec0c99",
          4082 => x"3d0d04da",
          4083 => x"3d0da93d",
          4084 => x"840551d2",
          4085 => x"f13f8253",
          4086 => x"a83dff84",
          4087 => x"0552a93d",
          4088 => x"51d5ee3f",
          4089 => x"828cec08",
          4090 => x"55828cec",
          4091 => x"0882d338",
          4092 => x"784da93d",
          4093 => x"08529d3d",
          4094 => x"705258cc",
          4095 => x"b83f828c",
          4096 => x"ec085582",
          4097 => x"8cec0882",
          4098 => x"b9380281",
          4099 => x"9b053381",
          4100 => x"a0065486",
          4101 => x"557382aa",
          4102 => x"38a053a4",
          4103 => x"3d0852a8",
          4104 => x"3dff8805",
          4105 => x"51ffb4ea",
          4106 => x"3fac5377",
          4107 => x"52923d70",
          4108 => x"5254ffb4",
          4109 => x"dd3faa3d",
          4110 => x"08527351",
          4111 => x"cbf73f82",
          4112 => x"8cec0855",
          4113 => x"828cec08",
          4114 => x"9538636f",
          4115 => x"2e098106",
          4116 => x"883865a2",
          4117 => x"3d082e92",
          4118 => x"38885581",
          4119 => x"e539828c",
          4120 => x"ec08842e",
          4121 => x"09810681",
          4122 => x"b8387351",
          4123 => x"c9b13f82",
          4124 => x"8cec0855",
          4125 => x"828cec08",
          4126 => x"81c83868",
          4127 => x"569353a8",
          4128 => x"3dff9505",
          4129 => x"528d1651",
          4130 => x"ffb4873f",
          4131 => x"02af0533",
          4132 => x"8b17348b",
          4133 => x"16337084",
          4134 => x"2a708106",
          4135 => x"51555573",
          4136 => x"893874a0",
          4137 => x"0754738b",
          4138 => x"17347854",
          4139 => x"810b8315",
          4140 => x"348b1633",
          4141 => x"70842a70",
          4142 => x"81065155",
          4143 => x"5573802e",
          4144 => x"80e5386e",
          4145 => x"642e80df",
          4146 => x"38755278",
          4147 => x"51c6be3f",
          4148 => x"828cec08",
          4149 => x"527851ff",
          4150 => x"b7bb3f82",
          4151 => x"55828cec",
          4152 => x"08802e80",
          4153 => x"dd38828c",
          4154 => x"ec085278",
          4155 => x"51ffb5af",
          4156 => x"3f828cec",
          4157 => x"087980d4",
          4158 => x"11585855",
          4159 => x"828cec08",
          4160 => x"80c03881",
          4161 => x"16335473",
          4162 => x"ae2e0981",
          4163 => x"06993863",
          4164 => x"53755276",
          4165 => x"51c6af3f",
          4166 => x"7854810b",
          4167 => x"83153487",
          4168 => x"39828cec",
          4169 => x"089c3877",
          4170 => x"51c8ca3f",
          4171 => x"828cec08",
          4172 => x"55828cec",
          4173 => x"088c3878",
          4174 => x"51ffb5aa",
          4175 => x"3f828cec",
          4176 => x"08557482",
          4177 => x"8cec0ca8",
          4178 => x"3d0d04ed",
          4179 => x"3d0d0280",
          4180 => x"db053302",
          4181 => x"840580df",
          4182 => x"05335757",
          4183 => x"8253953d",
          4184 => x"d0055296",
          4185 => x"3d51d2e9",
          4186 => x"3f828cec",
          4187 => x"0855828c",
          4188 => x"ec0880cf",
          4189 => x"38785a65",
          4190 => x"52953dd4",
          4191 => x"0551c9b5",
          4192 => x"3f828cec",
          4193 => x"0855828c",
          4194 => x"ec08b838",
          4195 => x"0280cf05",
          4196 => x"3381a006",
          4197 => x"54865573",
          4198 => x"aa3875a7",
          4199 => x"06617109",
          4200 => x"8b123371",
          4201 => x"067a7406",
          4202 => x"07515755",
          4203 => x"56748b15",
          4204 => x"34785481",
          4205 => x"0b831534",
          4206 => x"7851ffb4",
          4207 => x"a93f828c",
          4208 => x"ec085574",
          4209 => x"828cec0c",
          4210 => x"953d0d04",
          4211 => x"ef3d0d64",
          4212 => x"56825393",
          4213 => x"3dd00552",
          4214 => x"943d51d1",
          4215 => x"f43f828c",
          4216 => x"ec085582",
          4217 => x"8cec0880",
          4218 => x"cb387658",
          4219 => x"6352933d",
          4220 => x"d40551c8",
          4221 => x"c03f828c",
          4222 => x"ec085582",
          4223 => x"8cec08b4",
          4224 => x"380280c7",
          4225 => x"053381a0",
          4226 => x"06548655",
          4227 => x"73a63884",
          4228 => x"16228617",
          4229 => x"2271902b",
          4230 => x"07535496",
          4231 => x"1f51ffb0",
          4232 => x"c23f7654",
          4233 => x"810b8315",
          4234 => x"347651ff",
          4235 => x"b3b83f82",
          4236 => x"8cec0855",
          4237 => x"74828cec",
          4238 => x"0c933d0d",
          4239 => x"04ea3d0d",
          4240 => x"696b5c5a",
          4241 => x"8053983d",
          4242 => x"d0055299",
          4243 => x"3d51d181",
          4244 => x"3f828cec",
          4245 => x"08828cec",
          4246 => x"08307082",
          4247 => x"8cec0807",
          4248 => x"80255155",
          4249 => x"5779802e",
          4250 => x"81853881",
          4251 => x"70750655",
          4252 => x"5573802e",
          4253 => x"80f9387b",
          4254 => x"5d805f80",
          4255 => x"528d3d70",
          4256 => x"5254ffbe",
          4257 => x"a93f828c",
          4258 => x"ec085782",
          4259 => x"8cec0880",
          4260 => x"d1387452",
          4261 => x"7351c3dc",
          4262 => x"3f828cec",
          4263 => x"0857828c",
          4264 => x"ec08bf38",
          4265 => x"828cec08",
          4266 => x"828cec08",
          4267 => x"655b5956",
          4268 => x"78188119",
          4269 => x"7b185659",
          4270 => x"55743374",
          4271 => x"34811656",
          4272 => x"8a7827ec",
          4273 => x"388b5675",
          4274 => x"1a548074",
          4275 => x"3475802e",
          4276 => x"9e38ff16",
          4277 => x"701b7033",
          4278 => x"51555673",
          4279 => x"a02ee838",
          4280 => x"8e397684",
          4281 => x"2e098106",
          4282 => x"8638807a",
          4283 => x"34805776",
          4284 => x"30707807",
          4285 => x"80255154",
          4286 => x"7a802e80",
          4287 => x"c1387380",
          4288 => x"2ebc387b",
          4289 => x"a0110853",
          4290 => x"51ffb193",
          4291 => x"3f828cec",
          4292 => x"0857828c",
          4293 => x"ec08a738",
          4294 => x"7b703355",
          4295 => x"5580c356",
          4296 => x"73832e8b",
          4297 => x"3880e456",
          4298 => x"73842e83",
          4299 => x"38a75675",
          4300 => x"15b40551",
          4301 => x"ffade33f",
          4302 => x"828cec08",
          4303 => x"7b0c7682",
          4304 => x"8cec0c98",
          4305 => x"3d0d04e6",
          4306 => x"3d0d8253",
          4307 => x"9c3dffb8",
          4308 => x"05529d3d",
          4309 => x"51cefa3f",
          4310 => x"828cec08",
          4311 => x"828cec08",
          4312 => x"5654828c",
          4313 => x"ec088398",
          4314 => x"388b53a0",
          4315 => x"528b3d70",
          4316 => x"5259ffae",
          4317 => x"c03f736d",
          4318 => x"70337081",
          4319 => x"ff065257",
          4320 => x"55579f74",
          4321 => x"2781bc38",
          4322 => x"78587481",
          4323 => x"ff066d81",
          4324 => x"054e7052",
          4325 => x"55ffaf89",
          4326 => x"3f828cec",
          4327 => x"08802ea5",
          4328 => x"386c7033",
          4329 => x"70535754",
          4330 => x"ffaefd3f",
          4331 => x"828cec08",
          4332 => x"802e8d38",
          4333 => x"74882b76",
          4334 => x"076d8105",
          4335 => x"4e558639",
          4336 => x"828cec08",
          4337 => x"55ff9f15",
          4338 => x"7083ffff",
          4339 => x"06515473",
          4340 => x"99268a38",
          4341 => x"e0157083",
          4342 => x"ffff0656",
          4343 => x"5480ff75",
          4344 => x"27873881",
          4345 => x"fbbc1533",
          4346 => x"5574802e",
          4347 => x"a3387452",
          4348 => x"81fdbc51",
          4349 => x"ffae893f",
          4350 => x"828cec08",
          4351 => x"933881ff",
          4352 => x"75278838",
          4353 => x"76892688",
          4354 => x"388b398a",
          4355 => x"77278638",
          4356 => x"865581ec",
          4357 => x"3981ff75",
          4358 => x"278f3874",
          4359 => x"882a5473",
          4360 => x"78708105",
          4361 => x"5a348117",
          4362 => x"57747870",
          4363 => x"81055a34",
          4364 => x"81176d70",
          4365 => x"337081ff",
          4366 => x"06525755",
          4367 => x"57739f26",
          4368 => x"fec8388b",
          4369 => x"3d335486",
          4370 => x"557381e5",
          4371 => x"2e81b138",
          4372 => x"76802e99",
          4373 => x"3802a705",
          4374 => x"55761570",
          4375 => x"33515473",
          4376 => x"a02e0981",
          4377 => x"068738ff",
          4378 => x"175776ed",
          4379 => x"38794180",
          4380 => x"43805291",
          4381 => x"3d705255",
          4382 => x"ffbab33f",
          4383 => x"828cec08",
          4384 => x"54828cec",
          4385 => x"0880f738",
          4386 => x"81527451",
          4387 => x"ffbfe53f",
          4388 => x"828cec08",
          4389 => x"54828cec",
          4390 => x"088d3876",
          4391 => x"80c43867",
          4392 => x"54e57434",
          4393 => x"80c63982",
          4394 => x"8cec0884",
          4395 => x"2e098106",
          4396 => x"80cc3880",
          4397 => x"5476742e",
          4398 => x"80c43881",
          4399 => x"527451ff",
          4400 => x"bdb03f82",
          4401 => x"8cec0854",
          4402 => x"828cec08",
          4403 => x"b138a053",
          4404 => x"828cec08",
          4405 => x"526751ff",
          4406 => x"abdb3f67",
          4407 => x"54880b8b",
          4408 => x"15348b53",
          4409 => x"78526751",
          4410 => x"ffaba73f",
          4411 => x"7954810b",
          4412 => x"83153479",
          4413 => x"51ffadee",
          4414 => x"3f828cec",
          4415 => x"08547355",
          4416 => x"74828cec",
          4417 => x"0c9c3d0d",
          4418 => x"04f23d0d",
          4419 => x"60620288",
          4420 => x"0580cb05",
          4421 => x"33933dfc",
          4422 => x"05557254",
          4423 => x"405e5ad2",
          4424 => x"da3f828c",
          4425 => x"ec085882",
          4426 => x"8cec0882",
          4427 => x"bd38911a",
          4428 => x"33587782",
          4429 => x"b5387c80",
          4430 => x"2e97388c",
          4431 => x"1a085978",
          4432 => x"9038901a",
          4433 => x"3370812a",
          4434 => x"70810651",
          4435 => x"55557390",
          4436 => x"38875482",
          4437 => x"97398258",
          4438 => x"82903981",
          4439 => x"58828b39",
          4440 => x"7e8a1122",
          4441 => x"70892b70",
          4442 => x"557f5456",
          4443 => x"5656feff",
          4444 => x"c53fff14",
          4445 => x"7d067030",
          4446 => x"7072079f",
          4447 => x"2a828cec",
          4448 => x"08058c19",
          4449 => x"087c405a",
          4450 => x"5d555581",
          4451 => x"77278838",
          4452 => x"98160877",
          4453 => x"26833882",
          4454 => x"57767756",
          4455 => x"59805674",
          4456 => x"527951ff",
          4457 => x"ae993f81",
          4458 => x"157f5555",
          4459 => x"98140875",
          4460 => x"26833882",
          4461 => x"55828cec",
          4462 => x"08812eff",
          4463 => x"9938828c",
          4464 => x"ec08ff2e",
          4465 => x"ff953882",
          4466 => x"8cec088e",
          4467 => x"38811656",
          4468 => x"757b2e09",
          4469 => x"81068738",
          4470 => x"93397459",
          4471 => x"80567477",
          4472 => x"2e098106",
          4473 => x"ffb93887",
          4474 => x"5880ff39",
          4475 => x"7d802eba",
          4476 => x"38787b55",
          4477 => x"557a802e",
          4478 => x"b4388115",
          4479 => x"5673812e",
          4480 => x"09810683",
          4481 => x"38ff5675",
          4482 => x"5374527e",
          4483 => x"51ffafa8",
          4484 => x"3f828cec",
          4485 => x"0858828c",
          4486 => x"ec0880ce",
          4487 => x"38748116",
          4488 => x"ff165656",
          4489 => x"5c73d338",
          4490 => x"8439ff19",
          4491 => x"5c7e7c8c",
          4492 => x"120c557d",
          4493 => x"802eb338",
          4494 => x"78881b0c",
          4495 => x"7c8c1b0c",
          4496 => x"901a3380",
          4497 => x"c0075473",
          4498 => x"901b3498",
          4499 => x"1508fe05",
          4500 => x"90160857",
          4501 => x"54757426",
          4502 => x"9138757b",
          4503 => x"3190160c",
          4504 => x"84153381",
          4505 => x"07547384",
          4506 => x"16347754",
          4507 => x"73828cec",
          4508 => x"0c903d0d",
          4509 => x"04e93d0d",
          4510 => x"6b6d0288",
          4511 => x"0580eb05",
          4512 => x"339d3d54",
          4513 => x"5a5c59c5",
          4514 => x"bd3f8b56",
          4515 => x"800b828c",
          4516 => x"ec08248b",
          4517 => x"f838828c",
          4518 => x"ec088429",
          4519 => x"828d8805",
          4520 => x"70085155",
          4521 => x"74802e84",
          4522 => x"38807534",
          4523 => x"828cec08",
          4524 => x"81ff065f",
          4525 => x"81527e51",
          4526 => x"ffa0d03f",
          4527 => x"828cec08",
          4528 => x"81ff0670",
          4529 => x"81065657",
          4530 => x"8356748b",
          4531 => x"c0387682",
          4532 => x"2a708106",
          4533 => x"51558a56",
          4534 => x"748bb238",
          4535 => x"993dfc05",
          4536 => x"5383527e",
          4537 => x"51ffa4f0",
          4538 => x"3f828cec",
          4539 => x"08993867",
          4540 => x"5574802e",
          4541 => x"92387482",
          4542 => x"8080268b",
          4543 => x"38ff1575",
          4544 => x"06557480",
          4545 => x"2e833881",
          4546 => x"4878802e",
          4547 => x"87388480",
          4548 => x"79269238",
          4549 => x"7881800a",
          4550 => x"268b38ff",
          4551 => x"19790655",
          4552 => x"74802e86",
          4553 => x"3893568a",
          4554 => x"e4397889",
          4555 => x"2a6e892a",
          4556 => x"70892b77",
          4557 => x"59484359",
          4558 => x"7a833881",
          4559 => x"56613070",
          4560 => x"80257707",
          4561 => x"51559156",
          4562 => x"748ac238",
          4563 => x"993df805",
          4564 => x"5381527e",
          4565 => x"51ffa480",
          4566 => x"3f815682",
          4567 => x"8cec088a",
          4568 => x"ac387783",
          4569 => x"2a707706",
          4570 => x"828cec08",
          4571 => x"43564574",
          4572 => x"8338bf41",
          4573 => x"66558e56",
          4574 => x"6075268a",
          4575 => x"90387461",
          4576 => x"31704855",
          4577 => x"80ff7527",
          4578 => x"8a833893",
          4579 => x"56788180",
          4580 => x"2689fa38",
          4581 => x"77812a70",
          4582 => x"81065643",
          4583 => x"74802e95",
          4584 => x"38778706",
          4585 => x"5574822e",
          4586 => x"838d3877",
          4587 => x"81065574",
          4588 => x"802e8383",
          4589 => x"38778106",
          4590 => x"55935682",
          4591 => x"5e74802e",
          4592 => x"89cb3878",
          4593 => x"5a7d832e",
          4594 => x"09810680",
          4595 => x"e13878ae",
          4596 => x"3866912a",
          4597 => x"57810b81",
          4598 => x"fde02256",
          4599 => x"5a74802e",
          4600 => x"9d387477",
          4601 => x"26983881",
          4602 => x"fde05679",
          4603 => x"10821770",
          4604 => x"2257575a",
          4605 => x"74802e86",
          4606 => x"38767527",
          4607 => x"ee387952",
          4608 => x"6651fefa",
          4609 => x"b13f828c",
          4610 => x"ec088429",
          4611 => x"84870570",
          4612 => x"892a5e55",
          4613 => x"a05c800b",
          4614 => x"828cec08",
          4615 => x"fc808a05",
          4616 => x"5644fdff",
          4617 => x"f00a7527",
          4618 => x"80ec3888",
          4619 => x"d33978ae",
          4620 => x"38668c2a",
          4621 => x"57810b81",
          4622 => x"fdd02256",
          4623 => x"5a74802e",
          4624 => x"9d387477",
          4625 => x"26983881",
          4626 => x"fdd05679",
          4627 => x"10821770",
          4628 => x"2257575a",
          4629 => x"74802e86",
          4630 => x"38767527",
          4631 => x"ee387952",
          4632 => x"6651fef9",
          4633 => x"d13f828c",
          4634 => x"ec081084",
          4635 => x"0557828c",
          4636 => x"ec089ff5",
          4637 => x"26963881",
          4638 => x"0b828cec",
          4639 => x"0810828c",
          4640 => x"ec080571",
          4641 => x"11722a83",
          4642 => x"0559565e",
          4643 => x"83ff1789",
          4644 => x"2a5d815c",
          4645 => x"a044601c",
          4646 => x"7d116505",
          4647 => x"697012ff",
          4648 => x"05713070",
          4649 => x"72067431",
          4650 => x"5c525957",
          4651 => x"59407d83",
          4652 => x"2e098106",
          4653 => x"8938761c",
          4654 => x"6018415c",
          4655 => x"8439761d",
          4656 => x"5d799029",
          4657 => x"18706231",
          4658 => x"68585155",
          4659 => x"74762687",
          4660 => x"af38757c",
          4661 => x"317d317a",
          4662 => x"53706531",
          4663 => x"5255fef8",
          4664 => x"d53f828c",
          4665 => x"ec08587d",
          4666 => x"832e0981",
          4667 => x"069b3882",
          4668 => x"8cec0883",
          4669 => x"fff52680",
          4670 => x"dd387887",
          4671 => x"83387981",
          4672 => x"2a5978fd",
          4673 => x"be3886f8",
          4674 => x"397d822e",
          4675 => x"09810680",
          4676 => x"c53883ff",
          4677 => x"f50b828c",
          4678 => x"ec0827a0",
          4679 => x"38788f38",
          4680 => x"791a5574",
          4681 => x"80c02686",
          4682 => x"387459fd",
          4683 => x"96396281",
          4684 => x"06557480",
          4685 => x"2e8f3883",
          4686 => x"5efd8839",
          4687 => x"828cec08",
          4688 => x"9ff52692",
          4689 => x"387886b8",
          4690 => x"38791a59",
          4691 => x"81807927",
          4692 => x"fcf13886",
          4693 => x"ab398055",
          4694 => x"7d812e09",
          4695 => x"81068338",
          4696 => x"7d559ff5",
          4697 => x"78278b38",
          4698 => x"74810655",
          4699 => x"8e567486",
          4700 => x"9c388480",
          4701 => x"5380527a",
          4702 => x"51ffa2b9",
          4703 => x"3f8b5381",
          4704 => x"fbf8527a",
          4705 => x"51ffa28a",
          4706 => x"3f848052",
          4707 => x"8b1b51ff",
          4708 => x"a1b33f79",
          4709 => x"8d1c347b",
          4710 => x"83ffff06",
          4711 => x"528e1b51",
          4712 => x"ffa1a23f",
          4713 => x"810b901c",
          4714 => x"347d8332",
          4715 => x"70307096",
          4716 => x"2a848006",
          4717 => x"54515591",
          4718 => x"1b51ffa1",
          4719 => x"883f6655",
          4720 => x"7483ffff",
          4721 => x"26903874",
          4722 => x"83ffff06",
          4723 => x"52931b51",
          4724 => x"ffa0f23f",
          4725 => x"8a397452",
          4726 => x"a01b51ff",
          4727 => x"a1853ff8",
          4728 => x"0b951c34",
          4729 => x"bf52981b",
          4730 => x"51ffa0d9",
          4731 => x"3f81ff52",
          4732 => x"9a1b51ff",
          4733 => x"a0cf3f60",
          4734 => x"529c1b51",
          4735 => x"ffa0e43f",
          4736 => x"7d832e09",
          4737 => x"810680cb",
          4738 => x"388288b2",
          4739 => x"0a5280c3",
          4740 => x"1b51ffa0",
          4741 => x"ce3f7c52",
          4742 => x"a41b51ff",
          4743 => x"a0c53f82",
          4744 => x"52ac1b51",
          4745 => x"ffa0bc3f",
          4746 => x"8152b01b",
          4747 => x"51ffa095",
          4748 => x"3f8652b2",
          4749 => x"1b51ffa0",
          4750 => x"8c3fff80",
          4751 => x"0b80c01c",
          4752 => x"34a90b80",
          4753 => x"c21c3493",
          4754 => x"5381fc84",
          4755 => x"5280c71b",
          4756 => x"51ae3982",
          4757 => x"88b20a52",
          4758 => x"a71b51ff",
          4759 => x"a0853f7c",
          4760 => x"83ffff06",
          4761 => x"52961b51",
          4762 => x"ff9fda3f",
          4763 => x"ff800ba4",
          4764 => x"1c34a90b",
          4765 => x"a61c3493",
          4766 => x"5381fc98",
          4767 => x"52ab1b51",
          4768 => x"ffa08f3f",
          4769 => x"82d4d552",
          4770 => x"83fe1b70",
          4771 => x"5259ff9f",
          4772 => x"b43f8154",
          4773 => x"60537a52",
          4774 => x"7e51ff9b",
          4775 => x"d73f8156",
          4776 => x"828cec08",
          4777 => x"83e7387d",
          4778 => x"832e0981",
          4779 => x"0680ee38",
          4780 => x"75546086",
          4781 => x"05537a52",
          4782 => x"7e51ff9b",
          4783 => x"b73f8480",
          4784 => x"5380527a",
          4785 => x"51ff9fed",
          4786 => x"3f848b85",
          4787 => x"a4d2527a",
          4788 => x"51ff9f8f",
          4789 => x"3f868a85",
          4790 => x"e4f25283",
          4791 => x"e41b51ff",
          4792 => x"9f813fff",
          4793 => x"185283e8",
          4794 => x"1b51ff9e",
          4795 => x"f63f8252",
          4796 => x"83ec1b51",
          4797 => x"ff9eec3f",
          4798 => x"82d4d552",
          4799 => x"7851ff9e",
          4800 => x"c43f7554",
          4801 => x"60870553",
          4802 => x"7a527e51",
          4803 => x"ff9ae53f",
          4804 => x"75546016",
          4805 => x"537a527e",
          4806 => x"51ff9ad8",
          4807 => x"3f655380",
          4808 => x"527a51ff",
          4809 => x"9f8f3f7f",
          4810 => x"5680587d",
          4811 => x"832e0981",
          4812 => x"069a38f8",
          4813 => x"527a51ff",
          4814 => x"9ea93fff",
          4815 => x"52841b51",
          4816 => x"ff9ea03f",
          4817 => x"f00a5288",
          4818 => x"1b519139",
          4819 => x"87fffff8",
          4820 => x"557d812e",
          4821 => x"8338f855",
          4822 => x"74527a51",
          4823 => x"ff9e843f",
          4824 => x"7c556157",
          4825 => x"74622683",
          4826 => x"38745776",
          4827 => x"5475537a",
          4828 => x"527e51ff",
          4829 => x"99fe3f82",
          4830 => x"8cec0882",
          4831 => x"87388480",
          4832 => x"53828cec",
          4833 => x"08527a51",
          4834 => x"ff9eaa3f",
          4835 => x"76167578",
          4836 => x"31565674",
          4837 => x"cd388118",
          4838 => x"5877802e",
          4839 => x"ff8d3879",
          4840 => x"557d832e",
          4841 => x"83386355",
          4842 => x"61577462",
          4843 => x"26833874",
          4844 => x"57765475",
          4845 => x"537a527e",
          4846 => x"51ff99b8",
          4847 => x"3f828cec",
          4848 => x"0881c138",
          4849 => x"76167578",
          4850 => x"31565674",
          4851 => x"db388c56",
          4852 => x"7d832e93",
          4853 => x"38865666",
          4854 => x"83ffff26",
          4855 => x"8a388456",
          4856 => x"7d822e83",
          4857 => x"38815664",
          4858 => x"81065877",
          4859 => x"80fe3884",
          4860 => x"80537752",
          4861 => x"7a51ff9d",
          4862 => x"bc3f82d4",
          4863 => x"d5527851",
          4864 => x"ff9cc23f",
          4865 => x"83be1b55",
          4866 => x"77753481",
          4867 => x"0b811634",
          4868 => x"810b8216",
          4869 => x"34778316",
          4870 => x"34758416",
          4871 => x"34606705",
          4872 => x"5680fdc1",
          4873 => x"527551fe",
          4874 => x"f28c3ffe",
          4875 => x"0b851634",
          4876 => x"828cec08",
          4877 => x"822abf07",
          4878 => x"56758616",
          4879 => x"34828cec",
          4880 => x"08871634",
          4881 => x"605283c6",
          4882 => x"1b51ff9c",
          4883 => x"963f6652",
          4884 => x"83ca1b51",
          4885 => x"ff9c8c3f",
          4886 => x"81547753",
          4887 => x"7a527e51",
          4888 => x"ff98913f",
          4889 => x"8156828c",
          4890 => x"ec08a238",
          4891 => x"80538052",
          4892 => x"7e51ff99",
          4893 => x"e33f8156",
          4894 => x"828cec08",
          4895 => x"90388939",
          4896 => x"8e568a39",
          4897 => x"81568639",
          4898 => x"828cec08",
          4899 => x"5675828c",
          4900 => x"ec0c993d",
          4901 => x"0d04f53d",
          4902 => x"0d7d605b",
          4903 => x"59807960",
          4904 => x"ff055a57",
          4905 => x"57767825",
          4906 => x"b4388d3d",
          4907 => x"f8115555",
          4908 => x"8153fc15",
          4909 => x"527951c9",
          4910 => x"dc3f7a81",
          4911 => x"2e098106",
          4912 => x"9c388c3d",
          4913 => x"3355748d",
          4914 => x"2edb3874",
          4915 => x"76708105",
          4916 => x"58348117",
          4917 => x"57748a2e",
          4918 => x"098106c9",
          4919 => x"38807634",
          4920 => x"78557683",
          4921 => x"38765574",
          4922 => x"828cec0c",
          4923 => x"8d3d0d04",
          4924 => x"fa3d0d78",
          4925 => x"70087055",
          4926 => x"56577480",
          4927 => x"2e80ea38",
          4928 => x"8e397477",
          4929 => x"0c851433",
          4930 => x"5380de39",
          4931 => x"81155580",
          4932 => x"75335556",
          4933 => x"73a02e83",
          4934 => x"38815673",
          4935 => x"30709f2a",
          4936 => x"77065153",
          4937 => x"72e63873",
          4938 => x"a02e0981",
          4939 => x"06883872",
          4940 => x"75708105",
          4941 => x"57347256",
          4942 => x"75902982",
          4943 => x"89fc0577",
          4944 => x"08537008",
          4945 => x"5254fef3",
          4946 => x"f63f828c",
          4947 => x"ec088b38",
          4948 => x"84143353",
          4949 => x"72812eff",
          4950 => x"a9388116",
          4951 => x"7081ff06",
          4952 => x"57539676",
          4953 => x"27d238ff",
          4954 => x"5372828c",
          4955 => x"ec0c883d",
          4956 => x"0d04ff3d",
          4957 => x"0d735271",
          4958 => x"9326818e",
          4959 => x"38718429",
          4960 => x"81f59c05",
          4961 => x"52710804",
          4962 => x"81ff8851",
          4963 => x"81803981",
          4964 => x"ff945180",
          4965 => x"f93981ff",
          4966 => x"a85180f2",
          4967 => x"3981ffbc",
          4968 => x"5180eb39",
          4969 => x"81ffcc51",
          4970 => x"80e43981",
          4971 => x"ffdc5180",
          4972 => x"dd3981ff",
          4973 => x"f05180d6",
          4974 => x"39828080",
          4975 => x"5180cf39",
          4976 => x"82809851",
          4977 => x"80c83982",
          4978 => x"80b05180",
          4979 => x"c1398280",
          4980 => x"c851bb39",
          4981 => x"8280e451",
          4982 => x"b5398280",
          4983 => x"f851af39",
          4984 => x"8281a451",
          4985 => x"a9398281",
          4986 => x"b851a339",
          4987 => x"8281d851",
          4988 => x"9d398281",
          4989 => x"ec519739",
          4990 => x"82828451",
          4991 => x"91398282",
          4992 => x"9c518b39",
          4993 => x"8282b451",
          4994 => x"85398282",
          4995 => x"c051ff86",
          4996 => x"9f3f833d",
          4997 => x"0d04fb3d",
          4998 => x"0d777956",
          4999 => x"567487e7",
          5000 => x"268a3874",
          5001 => x"527587e8",
          5002 => x"29519139",
          5003 => x"87e85274",
          5004 => x"51feee82",
          5005 => x"3f828cec",
          5006 => x"08527551",
          5007 => x"feedf73f",
          5008 => x"828cec08",
          5009 => x"54795375",
          5010 => x"528282d0",
          5011 => x"51ff8bc4",
          5012 => x"3f873d0d",
          5013 => x"04ec3d0d",
          5014 => x"66028405",
          5015 => x"80e30533",
          5016 => x"5b578068",
          5017 => x"7830707a",
          5018 => x"07732551",
          5019 => x"57595978",
          5020 => x"567787ff",
          5021 => x"26833881",
          5022 => x"56747607",
          5023 => x"7081ff06",
          5024 => x"51559356",
          5025 => x"7480ff38",
          5026 => x"81537652",
          5027 => x"8c3d7052",
          5028 => x"56c19d3f",
          5029 => x"828cec08",
          5030 => x"57828cec",
          5031 => x"08b83882",
          5032 => x"8cec0887",
          5033 => x"c098880c",
          5034 => x"828cec08",
          5035 => x"59963dd4",
          5036 => x"05548480",
          5037 => x"53775275",
          5038 => x"51c5da3f",
          5039 => x"828cec08",
          5040 => x"57828cec",
          5041 => x"0890387a",
          5042 => x"5574802e",
          5043 => x"89387419",
          5044 => x"75195959",
          5045 => x"d839963d",
          5046 => x"d80551cd",
          5047 => x"c43f7630",
          5048 => x"70780780",
          5049 => x"257b3070",
          5050 => x"9f2a7206",
          5051 => x"51575156",
          5052 => x"74802e90",
          5053 => x"388282f4",
          5054 => x"5387c098",
          5055 => x"88085278",
          5056 => x"51fe933f",
          5057 => x"76567582",
          5058 => x"8cec0c96",
          5059 => x"3d0d04f9",
          5060 => x"3d0d7b02",
          5061 => x"8405b305",
          5062 => x"335758ff",
          5063 => x"5780537a",
          5064 => x"527951fe",
          5065 => x"b03f828c",
          5066 => x"ec08a438",
          5067 => x"75802e88",
          5068 => x"3875812e",
          5069 => x"98389839",
          5070 => x"60557f54",
          5071 => x"828cec53",
          5072 => x"7e527d51",
          5073 => x"772d828c",
          5074 => x"ec085783",
          5075 => x"39770476",
          5076 => x"828cec0c",
          5077 => x"893d0d04",
          5078 => x"f33d0d7f",
          5079 => x"6163028c",
          5080 => x"0580cf05",
          5081 => x"33737315",
          5082 => x"68415f5c",
          5083 => x"5c5e5e5e",
          5084 => x"7a528282",
          5085 => x"fc51ff89",
          5086 => x"9b3f8283",
          5087 => x"8451ff83",
          5088 => x"af3f8055",
          5089 => x"74792780",
          5090 => x"fc387b90",
          5091 => x"2e89387b",
          5092 => x"a02ea738",
          5093 => x"80c63974",
          5094 => x"1853727a",
          5095 => x"278e3872",
          5096 => x"22528283",
          5097 => x"8851ff88",
          5098 => x"eb3f8939",
          5099 => x"82839451",
          5100 => x"ff82fd3f",
          5101 => x"82155580",
          5102 => x"c3397418",
          5103 => x"53727a27",
          5104 => x"8e387208",
          5105 => x"528282fc",
          5106 => x"51ff88c8",
          5107 => x"3f893982",
          5108 => x"839051ff",
          5109 => x"82da3f84",
          5110 => x"1555a139",
          5111 => x"74185372",
          5112 => x"7a278e38",
          5113 => x"72335282",
          5114 => x"839c51ff",
          5115 => x"88a63f89",
          5116 => x"398283a4",
          5117 => x"51ff82b8",
          5118 => x"3f811555",
          5119 => x"a051ff81",
          5120 => x"d23fff80",
          5121 => x"398283a8",
          5122 => x"51ff82a4",
          5123 => x"3f805574",
          5124 => x"7927bc38",
          5125 => x"74187033",
          5126 => x"55538056",
          5127 => x"727a2783",
          5128 => x"38815680",
          5129 => x"539f7427",
          5130 => x"83388153",
          5131 => x"75730670",
          5132 => x"81ff0651",
          5133 => x"5372802e",
          5134 => x"8b387380",
          5135 => x"fe268538",
          5136 => x"73518339",
          5137 => x"a051ff81",
          5138 => x"8a3f8115",
          5139 => x"55c13982",
          5140 => x"83ac51ff",
          5141 => x"81da3f78",
          5142 => x"18791c5c",
          5143 => x"58fef6dc",
          5144 => x"3f828cec",
          5145 => x"08982b70",
          5146 => x"982c5157",
          5147 => x"76a02e09",
          5148 => x"8106ab38",
          5149 => x"fef6c53f",
          5150 => x"828cec08",
          5151 => x"982b7098",
          5152 => x"2c70a032",
          5153 => x"7030729b",
          5154 => x"32703070",
          5155 => x"72077375",
          5156 => x"07065158",
          5157 => x"58595751",
          5158 => x"57807324",
          5159 => x"d738769b",
          5160 => x"2e098106",
          5161 => x"85388053",
          5162 => x"8c397c1e",
          5163 => x"53727826",
          5164 => x"fdbe38ff",
          5165 => x"5372828c",
          5166 => x"ec0c8f3d",
          5167 => x"0d04fc3d",
          5168 => x"0d029b05",
          5169 => x"338283b0",
          5170 => x"538283b4",
          5171 => x"5255ff86",
          5172 => x"c33f8289",
          5173 => x"cc2251fe",
          5174 => x"ff9d3f82",
          5175 => x"83c05482",
          5176 => x"83cc5382",
          5177 => x"89cd3352",
          5178 => x"8283d451",
          5179 => x"ff86a53f",
          5180 => x"74802e85",
          5181 => x"38fefae8",
          5182 => x"3f863d0d",
          5183 => x"04fe3d0d",
          5184 => x"87c09680",
          5185 => x"0853feff",
          5186 => x"b83f8151",
          5187 => x"fef1c13f",
          5188 => x"8283f051",
          5189 => x"fef3b93f",
          5190 => x"8051fef1",
          5191 => x"b33f7281",
          5192 => x"2a708106",
          5193 => x"51527180",
          5194 => x"2e953881",
          5195 => x"51fef1a0",
          5196 => x"3f828488",
          5197 => x"51fef398",
          5198 => x"3f8051fe",
          5199 => x"f1923f72",
          5200 => x"822a7081",
          5201 => x"06515271",
          5202 => x"802e9538",
          5203 => x"8151fef0",
          5204 => x"ff3f8284",
          5205 => x"9c51fef2",
          5206 => x"f73f8051",
          5207 => x"fef0f13f",
          5208 => x"72832a70",
          5209 => x"81065152",
          5210 => x"71802e95",
          5211 => x"388151fe",
          5212 => x"f0de3f82",
          5213 => x"84ac51fe",
          5214 => x"f2d63f80",
          5215 => x"51fef0d0",
          5216 => x"3f72842a",
          5217 => x"70810651",
          5218 => x"5271802e",
          5219 => x"95388151",
          5220 => x"fef0bd3f",
          5221 => x"8284c051",
          5222 => x"fef2b53f",
          5223 => x"8051fef0",
          5224 => x"af3f7285",
          5225 => x"2a708106",
          5226 => x"51527180",
          5227 => x"2e953881",
          5228 => x"51fef09c",
          5229 => x"3f8284d4",
          5230 => x"51fef294",
          5231 => x"3f8051fe",
          5232 => x"f08e3f72",
          5233 => x"862a7081",
          5234 => x"06515271",
          5235 => x"802e9538",
          5236 => x"8151feef",
          5237 => x"fb3f8284",
          5238 => x"e851fef1",
          5239 => x"f33f8051",
          5240 => x"feefed3f",
          5241 => x"72872a70",
          5242 => x"81065152",
          5243 => x"71802e95",
          5244 => x"388151fe",
          5245 => x"efda3f82",
          5246 => x"84fc51fe",
          5247 => x"f1d23f80",
          5248 => x"51feefcc",
          5249 => x"3f72882a",
          5250 => x"70810651",
          5251 => x"5271802e",
          5252 => x"95388151",
          5253 => x"feefb93f",
          5254 => x"82859051",
          5255 => x"fef1b13f",
          5256 => x"8051feef",
          5257 => x"ab3ffefd",
          5258 => x"a03f843d",
          5259 => x"0d04fb3d",
          5260 => x"0d777970",
          5261 => x"55565680",
          5262 => x"527551fe",
          5263 => x"e8f03f82",
          5264 => x"89f83354",
          5265 => x"73a73881",
          5266 => x"538285d0",
          5267 => x"5282a3f0",
          5268 => x"51ffb9dc",
          5269 => x"3f828cec",
          5270 => x"08307082",
          5271 => x"8cec0807",
          5272 => x"80258271",
          5273 => x"31515154",
          5274 => x"738289f8",
          5275 => x"348289f8",
          5276 => x"33547381",
          5277 => x"2e098106",
          5278 => x"ac3882a3",
          5279 => x"f0537452",
          5280 => x"7551f492",
          5281 => x"3f828cec",
          5282 => x"08802e8c",
          5283 => x"38828cec",
          5284 => x"0851fefd",
          5285 => x"9b3f8e39",
          5286 => x"82a3f051",
          5287 => x"c6833f82",
          5288 => x"0b8289f8",
          5289 => x"348289f8",
          5290 => x"33547382",
          5291 => x"2e098106",
          5292 => x"89387452",
          5293 => x"7551ff83",
          5294 => x"b53f800b",
          5295 => x"828cec0c",
          5296 => x"873d0d04",
          5297 => x"ce3d0d80",
          5298 => x"707182a3",
          5299 => x"ec0c5f5d",
          5300 => x"81527c51",
          5301 => x"ff88b43f",
          5302 => x"828cec08",
          5303 => x"81ff0659",
          5304 => x"787d2e09",
          5305 => x"8106a238",
          5306 => x"8285e052",
          5307 => x"963d7052",
          5308 => x"59ff82b6",
          5309 => x"3f7c5378",
          5310 => x"52828e9c",
          5311 => x"51ffb7cf",
          5312 => x"3f828cec",
          5313 => x"087d2e88",
          5314 => x"388285e4",
          5315 => x"518dc139",
          5316 => x"81705f5d",
          5317 => x"82869c51",
          5318 => x"fefc953f",
          5319 => x"963d7046",
          5320 => x"5a80f852",
          5321 => x"7951fe86",
          5322 => x"3fb43dff",
          5323 => x"840551f3",
          5324 => x"bf3f828c",
          5325 => x"ec08902b",
          5326 => x"70902c51",
          5327 => x"597880c2",
          5328 => x"2e87b338",
          5329 => x"7880c224",
          5330 => x"b23878bd",
          5331 => x"2e81d538",
          5332 => x"78bd2490",
          5333 => x"3878802e",
          5334 => x"ffba3878",
          5335 => x"bc2e80da",
          5336 => x"388ae939",
          5337 => x"7880c02e",
          5338 => x"83a13878",
          5339 => x"80c02485",
          5340 => x"dd3878bf",
          5341 => x"2e829238",
          5342 => x"8ad23978",
          5343 => x"80f92e89",
          5344 => x"ea387880",
          5345 => x"f9249238",
          5346 => x"7880c32e",
          5347 => x"88983878",
          5348 => x"80f82e89",
          5349 => x"b1388ab4",
          5350 => x"39788183",
          5351 => x"2e8a9938",
          5352 => x"78818324",
          5353 => x"8b387881",
          5354 => x"822e89fd",
          5355 => x"388a9d39",
          5356 => x"7881852e",
          5357 => x"8a8f388a",
          5358 => x"9339b43d",
          5359 => x"ff801153",
          5360 => x"ff840551",
          5361 => x"ff82c23f",
          5362 => x"828cec08",
          5363 => x"802efec4",
          5364 => x"38b43dfe",
          5365 => x"fc1153ff",
          5366 => x"840551ff",
          5367 => x"82ab3f82",
          5368 => x"8cec0880",
          5369 => x"2efead38",
          5370 => x"b43dfef8",
          5371 => x"1153ff84",
          5372 => x"0551ff82",
          5373 => x"943f828c",
          5374 => x"ec088638",
          5375 => x"828cec08",
          5376 => x"428286a0",
          5377 => x"51fefaa8",
          5378 => x"3f63635c",
          5379 => x"5a797b27",
          5380 => x"81f23861",
          5381 => x"59787a70",
          5382 => x"84055c0c",
          5383 => x"7a7a26f5",
          5384 => x"3881e139",
          5385 => x"b43dff80",
          5386 => x"1153ff84",
          5387 => x"0551ff81",
          5388 => x"d83f828c",
          5389 => x"ec08802e",
          5390 => x"fdda38b4",
          5391 => x"3dfefc11",
          5392 => x"53ff8405",
          5393 => x"51ff81c1",
          5394 => x"3f828cec",
          5395 => x"08802efd",
          5396 => x"c338b43d",
          5397 => x"fef81153",
          5398 => x"ff840551",
          5399 => x"ff81aa3f",
          5400 => x"828cec08",
          5401 => x"802efdac",
          5402 => x"388286b0",
          5403 => x"51fef9c0",
          5404 => x"3f635a79",
          5405 => x"6327818c",
          5406 => x"38615979",
          5407 => x"7081055b",
          5408 => x"33793461",
          5409 => x"810542eb",
          5410 => x"39b43dff",
          5411 => x"801153ff",
          5412 => x"840551ff",
          5413 => x"80f33f82",
          5414 => x"8cec0880",
          5415 => x"2efcf538",
          5416 => x"b43dfefc",
          5417 => x"1153ff84",
          5418 => x"0551ff80",
          5419 => x"dc3f828c",
          5420 => x"ec08802e",
          5421 => x"fcde38b4",
          5422 => x"3dfef811",
          5423 => x"53ff8405",
          5424 => x"51ff80c5",
          5425 => x"3f828cec",
          5426 => x"08802efc",
          5427 => x"c7388286",
          5428 => x"bc51fef8",
          5429 => x"db3f635a",
          5430 => x"796327a8",
          5431 => x"38617033",
          5432 => x"7b335e5a",
          5433 => x"5b787c2e",
          5434 => x"92387855",
          5435 => x"7a547933",
          5436 => x"53795282",
          5437 => x"86cc51fe",
          5438 => x"fe9a3f81",
          5439 => x"1a628105",
          5440 => x"435ad539",
          5441 => x"8286e451",
          5442 => x"82bd39b4",
          5443 => x"3dff8011",
          5444 => x"53ff8405",
          5445 => x"51fefff1",
          5446 => x"3f828cec",
          5447 => x"0880df38",
          5448 => x"8289e033",
          5449 => x"5978802e",
          5450 => x"89388289",
          5451 => x"98084480",
          5452 => x"cd398289",
          5453 => x"e1335978",
          5454 => x"802e8838",
          5455 => x"8289a008",
          5456 => x"44bc3982",
          5457 => x"89e23359",
          5458 => x"78802e88",
          5459 => x"388289a8",
          5460 => x"0844ab39",
          5461 => x"8289e333",
          5462 => x"5978802e",
          5463 => x"88388289",
          5464 => x"b008449a",
          5465 => x"398289de",
          5466 => x"33597880",
          5467 => x"2e883882",
          5468 => x"89b80844",
          5469 => x"89398289",
          5470 => x"c808fc80",
          5471 => x"0544b43d",
          5472 => x"fefc1153",
          5473 => x"ff840551",
          5474 => x"fefefe3f",
          5475 => x"828cec08",
          5476 => x"80de3882",
          5477 => x"89e03359",
          5478 => x"78802e89",
          5479 => x"3882899c",
          5480 => x"084380cc",
          5481 => x"398289e1",
          5482 => x"33597880",
          5483 => x"2e883882",
          5484 => x"89a40843",
          5485 => x"bb398289",
          5486 => x"e2335978",
          5487 => x"802e8838",
          5488 => x"8289ac08",
          5489 => x"43aa3982",
          5490 => x"89e33359",
          5491 => x"78802e88",
          5492 => x"388289b4",
          5493 => x"08439939",
          5494 => x"8289de33",
          5495 => x"5978802e",
          5496 => x"88388289",
          5497 => x"bc084388",
          5498 => x"398289c8",
          5499 => x"08880543",
          5500 => x"b43dfef8",
          5501 => x"1153ff84",
          5502 => x"0551fefe",
          5503 => x"8c3f828c",
          5504 => x"ec08802e",
          5505 => x"a7388062",
          5506 => x"5c5c7a88",
          5507 => x"2e833881",
          5508 => x"5c7a9032",
          5509 => x"70307072",
          5510 => x"079f2a70",
          5511 => x"7f065151",
          5512 => x"5a5a7880",
          5513 => x"2e88387a",
          5514 => x"a02e8338",
          5515 => x"88428286",
          5516 => x"e851fef5",
          5517 => x"fb3fa055",
          5518 => x"63546153",
          5519 => x"62526351",
          5520 => x"f2963f82",
          5521 => x"86f851fe",
          5522 => x"f5e63ff9",
          5523 => x"c739b43d",
          5524 => x"ff801153",
          5525 => x"ff840551",
          5526 => x"fefdae3f",
          5527 => x"828cec08",
          5528 => x"802ef9b0",
          5529 => x"38b43dfe",
          5530 => x"fc1153ff",
          5531 => x"840551fe",
          5532 => x"fd973f82",
          5533 => x"8cec0880",
          5534 => x"2ea53863",
          5535 => x"590280cb",
          5536 => x"05337934",
          5537 => x"63810544",
          5538 => x"b43dfefc",
          5539 => x"1153ff84",
          5540 => x"0551fefc",
          5541 => x"f43f828c",
          5542 => x"ec08e038",
          5543 => x"f8f63963",
          5544 => x"70335452",
          5545 => x"82878451",
          5546 => x"fefae93f",
          5547 => x"80f85279",
          5548 => x"51fefbba",
          5549 => x"3f794579",
          5550 => x"335978ae",
          5551 => x"2ef8d538",
          5552 => x"9f7927a0",
          5553 => x"38b43dfe",
          5554 => x"fc1153ff",
          5555 => x"840551fe",
          5556 => x"fcb73f82",
          5557 => x"8cec0880",
          5558 => x"2e913863",
          5559 => x"590280cb",
          5560 => x"05337934",
          5561 => x"63810544",
          5562 => x"ffb53982",
          5563 => x"879051fe",
          5564 => x"f4be3fff",
          5565 => x"aa39b43d",
          5566 => x"fef41153",
          5567 => x"ff840551",
          5568 => x"fefdf83f",
          5569 => x"828cec08",
          5570 => x"802ef888",
          5571 => x"38b43dfe",
          5572 => x"f01153ff",
          5573 => x"840551fe",
          5574 => x"fde13f82",
          5575 => x"8cec0880",
          5576 => x"2ea63860",
          5577 => x"5902be05",
          5578 => x"22797082",
          5579 => x"055b2378",
          5580 => x"41b43dfe",
          5581 => x"f01153ff",
          5582 => x"840551fe",
          5583 => x"fdbd3f82",
          5584 => x"8cec08df",
          5585 => x"38f7cd39",
          5586 => x"60702254",
          5587 => x"52828798",
          5588 => x"51fef9c0",
          5589 => x"3f80f852",
          5590 => x"7951fefa",
          5591 => x"913f7945",
          5592 => x"79335978",
          5593 => x"ae2ef7ac",
          5594 => x"38789f26",
          5595 => x"87386082",
          5596 => x"0541d539",
          5597 => x"b43dfef0",
          5598 => x"1153ff84",
          5599 => x"0551fefc",
          5600 => x"fa3f828c",
          5601 => x"ec08802e",
          5602 => x"92386059",
          5603 => x"02be0522",
          5604 => x"79708205",
          5605 => x"5b237841",
          5606 => x"ffae3982",
          5607 => x"879051fe",
          5608 => x"f38e3fff",
          5609 => x"a339b43d",
          5610 => x"fef41153",
          5611 => x"ff840551",
          5612 => x"fefcc83f",
          5613 => x"828cec08",
          5614 => x"802ef6d8",
          5615 => x"38b43dfe",
          5616 => x"f01153ff",
          5617 => x"840551fe",
          5618 => x"fcb13f82",
          5619 => x"8cec0880",
          5620 => x"2ea13860",
          5621 => x"60710c59",
          5622 => x"60840541",
          5623 => x"b43dfef0",
          5624 => x"1153ff84",
          5625 => x"0551fefc",
          5626 => x"923f828c",
          5627 => x"ec08e438",
          5628 => x"f6a23960",
          5629 => x"70085452",
          5630 => x"8287a451",
          5631 => x"fef8953f",
          5632 => x"80f85279",
          5633 => x"51fef8e6",
          5634 => x"3f794579",
          5635 => x"335978ae",
          5636 => x"2ef68138",
          5637 => x"9f79279c",
          5638 => x"38b43dfe",
          5639 => x"f01153ff",
          5640 => x"840551fe",
          5641 => x"fbd53f82",
          5642 => x"8cec0880",
          5643 => x"2e8d3860",
          5644 => x"60710c59",
          5645 => x"60840541",
          5646 => x"ffb93982",
          5647 => x"879051fe",
          5648 => x"f1ee3fff",
          5649 => x"ae39b43d",
          5650 => x"ff801153",
          5651 => x"ff840551",
          5652 => x"fef9b63f",
          5653 => x"828cec08",
          5654 => x"802ef5b8",
          5655 => x"38635282",
          5656 => x"87b051fe",
          5657 => x"f7ae3f63",
          5658 => x"597804b4",
          5659 => x"3dff8011",
          5660 => x"53ff8405",
          5661 => x"51fef991",
          5662 => x"3f828cec",
          5663 => x"08802ef5",
          5664 => x"93386352",
          5665 => x"8287cc51",
          5666 => x"fef7893f",
          5667 => x"6359782d",
          5668 => x"828cec08",
          5669 => x"802ef4fc",
          5670 => x"38828cec",
          5671 => x"08528287",
          5672 => x"e851fef6",
          5673 => x"ef3ff4ec",
          5674 => x"39828884",
          5675 => x"51fef180",
          5676 => x"3ffed8e1",
          5677 => x"3ff4dd39",
          5678 => x"8288a051",
          5679 => x"fef0f13f",
          5680 => x"8059ffa5",
          5681 => x"39feeb98",
          5682 => x"3ff4c939",
          5683 => x"64703351",
          5684 => x"5978802e",
          5685 => x"f4be387d",
          5686 => x"7d065978",
          5687 => x"802e81d8",
          5688 => x"38b43dff",
          5689 => x"840551fe",
          5690 => x"de973f82",
          5691 => x"8cec085c",
          5692 => x"815b7a82",
          5693 => x"2eb2387a",
          5694 => x"82248938",
          5695 => x"7a812e8c",
          5696 => x"3880cd39",
          5697 => x"7a832eb0",
          5698 => x"3880c539",
          5699 => x"8288b456",
          5700 => x"7b558288",
          5701 => x"b8548053",
          5702 => x"8288bc52",
          5703 => x"b43dffb0",
          5704 => x"0551fef6",
          5705 => x"853fbb39",
          5706 => x"8288dc52",
          5707 => x"b43dffb0",
          5708 => x"0551fef5",
          5709 => x"f53fab39",
          5710 => x"7b558288",
          5711 => x"b8548053",
          5712 => x"8288cc52",
          5713 => x"b43dffb0",
          5714 => x"0551fef5",
          5715 => x"dd3f9339",
          5716 => x"7b548053",
          5717 => x"8288d852",
          5718 => x"b43dffb0",
          5719 => x"0551fef5",
          5720 => x"c93f8289",
          5721 => x"9858828d",
          5722 => x"a0578056",
          5723 => x"64811146",
          5724 => x"81055580",
          5725 => x"54838080",
          5726 => x"53838080",
          5727 => x"52b43dff",
          5728 => x"b00551eb",
          5729 => x"8a3f828c",
          5730 => x"ec08828c",
          5731 => x"ec080970",
          5732 => x"30707207",
          5733 => x"8025515b",
          5734 => x"5b5f805a",
          5735 => x"7a832683",
          5736 => x"38815a78",
          5737 => x"7a065978",
          5738 => x"802e8d38",
          5739 => x"811b7081",
          5740 => x"ff065c59",
          5741 => x"7afebb38",
          5742 => x"7d81327d",
          5743 => x"81320759",
          5744 => x"788a387e",
          5745 => x"ff2e0981",
          5746 => x"06f2c938",
          5747 => x"8288e051",
          5748 => x"fef4c13f",
          5749 => x"f2be39fc",
          5750 => x"3d0d800b",
          5751 => x"828da034",
          5752 => x"87c0948c",
          5753 => x"70085455",
          5754 => x"87848052",
          5755 => x"7251fed6",
          5756 => x"c53f828c",
          5757 => x"ec08902b",
          5758 => x"75085553",
          5759 => x"87848052",
          5760 => x"7351fed6",
          5761 => x"b13f7282",
          5762 => x"8cec0807",
          5763 => x"750c87c0",
          5764 => x"949c7008",
          5765 => x"54558784",
          5766 => x"80527251",
          5767 => x"fed6973f",
          5768 => x"828cec08",
          5769 => x"902b7508",
          5770 => x"55538784",
          5771 => x"80527351",
          5772 => x"fed6833f",
          5773 => x"72828cec",
          5774 => x"0807750c",
          5775 => x"8c80830b",
          5776 => x"87c09484",
          5777 => x"0c8c8083",
          5778 => x"0b87c094",
          5779 => x"940c80d3",
          5780 => x"ea0b828c",
          5781 => x"fc0c80d6",
          5782 => x"eb0b828d",
          5783 => x"800cfee3",
          5784 => x"b33ffeec",
          5785 => x"dc3f8288",
          5786 => x"f051feed",
          5787 => x"c33f8288",
          5788 => x"fc51feed",
          5789 => x"bb3f81e1",
          5790 => x"fd51feec",
          5791 => x"bf3f8151",
          5792 => x"ecbc3ff0",
          5793 => x"bf3f8004",
          5794 => x"00003093",
          5795 => x"00003099",
          5796 => x"0000309f",
          5797 => x"000030a5",
          5798 => x"000030ab",
          5799 => x"00006e04",
          5800 => x"00006d88",
          5801 => x"00006d8f",
          5802 => x"00006d96",
          5803 => x"00006d9d",
          5804 => x"00006da4",
          5805 => x"00006dab",
          5806 => x"00006db2",
          5807 => x"00006db9",
          5808 => x"00006dc0",
          5809 => x"00006dc7",
          5810 => x"00006dce",
          5811 => x"00006dd4",
          5812 => x"00006dda",
          5813 => x"00006de0",
          5814 => x"00006de6",
          5815 => x"00006dec",
          5816 => x"00006df2",
          5817 => x"00006df8",
          5818 => x"00006dfe",
          5819 => x"25642f25",
          5820 => x"642f2564",
          5821 => x"2025643a",
          5822 => x"25643a25",
          5823 => x"642e2564",
          5824 => x"25640a00",
          5825 => x"536f4320",
          5826 => x"436f6e66",
          5827 => x"69677572",
          5828 => x"6174696f",
          5829 => x"6e000000",
          5830 => x"20286672",
          5831 => x"6f6d2053",
          5832 => x"6f432063",
          5833 => x"6f6e6669",
          5834 => x"67290000",
          5835 => x"3a0a4465",
          5836 => x"76696365",
          5837 => x"7320696d",
          5838 => x"706c656d",
          5839 => x"656e7465",
          5840 => x"643a0a00",
          5841 => x"20202020",
          5842 => x"57422053",
          5843 => x"4452414d",
          5844 => x"20202825",
          5845 => x"3038583a",
          5846 => x"25303858",
          5847 => x"292e0a00",
          5848 => x"20202020",
          5849 => x"53445241",
          5850 => x"4d202020",
          5851 => x"20202825",
          5852 => x"3038583a",
          5853 => x"25303858",
          5854 => x"292e0a00",
          5855 => x"20202020",
          5856 => x"494e534e",
          5857 => x"20425241",
          5858 => x"4d202825",
          5859 => x"3038583a",
          5860 => x"25303858",
          5861 => x"292e0a00",
          5862 => x"20202020",
          5863 => x"4252414d",
          5864 => x"20202020",
          5865 => x"20202825",
          5866 => x"3038583a",
          5867 => x"25303858",
          5868 => x"292e0a00",
          5869 => x"20202020",
          5870 => x"52414d20",
          5871 => x"20202020",
          5872 => x"20202825",
          5873 => x"3038583a",
          5874 => x"25303858",
          5875 => x"292e0a00",
          5876 => x"20202020",
          5877 => x"53442043",
          5878 => x"41524420",
          5879 => x"20202844",
          5880 => x"65766963",
          5881 => x"6573203d",
          5882 => x"25303264",
          5883 => x"292e0a00",
          5884 => x"20202020",
          5885 => x"54494d45",
          5886 => x"52312020",
          5887 => x"20202854",
          5888 => x"696d6572",
          5889 => x"7320203d",
          5890 => x"25303264",
          5891 => x"292e0a00",
          5892 => x"20202020",
          5893 => x"494e5452",
          5894 => x"20435452",
          5895 => x"4c202843",
          5896 => x"68616e6e",
          5897 => x"656c733d",
          5898 => x"25303264",
          5899 => x"292e0a00",
          5900 => x"20202020",
          5901 => x"57495348",
          5902 => x"424f4e45",
          5903 => x"20425553",
          5904 => x"0a000000",
          5905 => x"20202020",
          5906 => x"57422049",
          5907 => x"32430a00",
          5908 => x"20202020",
          5909 => x"494f4354",
          5910 => x"4c0a0000",
          5911 => x"20202020",
          5912 => x"5053320a",
          5913 => x"00000000",
          5914 => x"20202020",
          5915 => x"5350490a",
          5916 => x"00000000",
          5917 => x"41646472",
          5918 => x"65737365",
          5919 => x"733a0a00",
          5920 => x"20202020",
          5921 => x"43505520",
          5922 => x"52657365",
          5923 => x"74205665",
          5924 => x"63746f72",
          5925 => x"20416464",
          5926 => x"72657373",
          5927 => x"203d2025",
          5928 => x"3038580a",
          5929 => x"00000000",
          5930 => x"20202020",
          5931 => x"43505520",
          5932 => x"4d656d6f",
          5933 => x"72792053",
          5934 => x"74617274",
          5935 => x"20416464",
          5936 => x"72657373",
          5937 => x"203d2025",
          5938 => x"3038580a",
          5939 => x"00000000",
          5940 => x"20202020",
          5941 => x"53746163",
          5942 => x"6b205374",
          5943 => x"61727420",
          5944 => x"41646472",
          5945 => x"65737320",
          5946 => x"20202020",
          5947 => x"203d2025",
          5948 => x"3038580a",
          5949 => x"00000000",
          5950 => x"4d697363",
          5951 => x"3a0a0000",
          5952 => x"20202020",
          5953 => x"5a505520",
          5954 => x"49642020",
          5955 => x"20202020",
          5956 => x"20202020",
          5957 => x"20202020",
          5958 => x"20202020",
          5959 => x"203d2025",
          5960 => x"3034580a",
          5961 => x"00000000",
          5962 => x"20202020",
          5963 => x"53797374",
          5964 => x"656d2043",
          5965 => x"6c6f636b",
          5966 => x"20467265",
          5967 => x"71202020",
          5968 => x"20202020",
          5969 => x"203d2025",
          5970 => x"642e2530",
          5971 => x"34644d48",
          5972 => x"7a0a0000",
          5973 => x"20202020",
          5974 => x"53445241",
          5975 => x"4d20436c",
          5976 => x"6f636b20",
          5977 => x"46726571",
          5978 => x"20202020",
          5979 => x"20202020",
          5980 => x"203d2025",
          5981 => x"642e2530",
          5982 => x"34644d48",
          5983 => x"7a0a0000",
          5984 => x"20202020",
          5985 => x"57697368",
          5986 => x"626f6e65",
          5987 => x"20534452",
          5988 => x"414d2043",
          5989 => x"6c6f636b",
          5990 => x"20467265",
          5991 => x"713d2025",
          5992 => x"642e2530",
          5993 => x"34644d48",
          5994 => x"7a0a0000",
          5995 => x"536d616c",
          5996 => x"6c000000",
          5997 => x"4d656469",
          5998 => x"756d0000",
          5999 => x"466c6578",
          6000 => x"00000000",
          6001 => x"45564f00",
          6002 => x"45564f6d",
          6003 => x"696e0000",
          6004 => x"556e6b6e",
          6005 => x"6f776e00",
          6006 => x"53440000",
          6007 => x"222a2b2c",
          6008 => x"3a3b3c3d",
          6009 => x"3e3f5b5d",
          6010 => x"7c7f0000",
          6011 => x"46415400",
          6012 => x"46415433",
          6013 => x"32000000",
          6014 => x"ebfe904d",
          6015 => x"53444f53",
          6016 => x"352e3000",
          6017 => x"4e4f204e",
          6018 => x"414d4520",
          6019 => x"20202046",
          6020 => x"41543332",
          6021 => x"20202000",
          6022 => x"4e4f204e",
          6023 => x"414d4520",
          6024 => x"20202046",
          6025 => x"41542020",
          6026 => x"20202000",
          6027 => x"00007dd8",
          6028 => x"00000000",
          6029 => x"00000000",
          6030 => x"00000000",
          6031 => x"809a4541",
          6032 => x"8e418f80",
          6033 => x"45454549",
          6034 => x"49498e8f",
          6035 => x"9092924f",
          6036 => x"994f5555",
          6037 => x"59999a9b",
          6038 => x"9c9d9e9f",
          6039 => x"41494f55",
          6040 => x"a5a5a6a7",
          6041 => x"a8a9aaab",
          6042 => x"acadaeaf",
          6043 => x"b0b1b2b3",
          6044 => x"b4b5b6b7",
          6045 => x"b8b9babb",
          6046 => x"bcbdbebf",
          6047 => x"c0c1c2c3",
          6048 => x"c4c5c6c7",
          6049 => x"c8c9cacb",
          6050 => x"cccdcecf",
          6051 => x"d0d1d2d3",
          6052 => x"d4d5d6d7",
          6053 => x"d8d9dadb",
          6054 => x"dcdddedf",
          6055 => x"e0e1e2e3",
          6056 => x"e4e5e6e7",
          6057 => x"e8e9eaeb",
          6058 => x"ecedeeef",
          6059 => x"f0f1f2f3",
          6060 => x"f4f5f6f7",
          6061 => x"f8f9fafb",
          6062 => x"fcfdfeff",
          6063 => x"2b2e2c3b",
          6064 => x"3d5b5d2f",
          6065 => x"5c222a3a",
          6066 => x"3c3e3f7c",
          6067 => x"7f000000",
          6068 => x"00010004",
          6069 => x"00100040",
          6070 => x"01000200",
          6071 => x"00000000",
          6072 => x"00010002",
          6073 => x"00040008",
          6074 => x"00100020",
          6075 => x"00000000",
          6076 => x"64696e69",
          6077 => x"74000000",
          6078 => x"64696f63",
          6079 => x"746c0000",
          6080 => x"66696e69",
          6081 => x"74000000",
          6082 => x"666c6f61",
          6083 => x"64000000",
          6084 => x"66657865",
          6085 => x"63000000",
          6086 => x"6d636c65",
          6087 => x"61720000",
          6088 => x"6d636f70",
          6089 => x"79000000",
          6090 => x"6d646966",
          6091 => x"66000000",
          6092 => x"6d64756d",
          6093 => x"70000000",
          6094 => x"6d656200",
          6095 => x"6d656800",
          6096 => x"6d657700",
          6097 => x"68696400",
          6098 => x"68696500",
          6099 => x"68666400",
          6100 => x"68666500",
          6101 => x"63616c6c",
          6102 => x"00000000",
          6103 => x"6a6d7000",
          6104 => x"72657374",
          6105 => x"61727400",
          6106 => x"72657365",
          6107 => x"74000000",
          6108 => x"696e666f",
          6109 => x"00000000",
          6110 => x"74657374",
          6111 => x"00000000",
          6112 => x"74626173",
          6113 => x"69630000",
          6114 => x"4469736b",
          6115 => x"20457272",
          6116 => x"6f720a00",
          6117 => x"496e7465",
          6118 => x"726e616c",
          6119 => x"20657272",
          6120 => x"6f722e0a",
          6121 => x"00000000",
          6122 => x"4469736b",
          6123 => x"206e6f74",
          6124 => x"20726561",
          6125 => x"64792e0a",
          6126 => x"00000000",
          6127 => x"4e6f2066",
          6128 => x"696c6520",
          6129 => x"666f756e",
          6130 => x"642e0a00",
          6131 => x"4e6f2070",
          6132 => x"61746820",
          6133 => x"666f756e",
          6134 => x"642e0a00",
          6135 => x"496e7661",
          6136 => x"6c696420",
          6137 => x"66696c65",
          6138 => x"6e616d65",
          6139 => x"2e0a0000",
          6140 => x"41636365",
          6141 => x"73732064",
          6142 => x"656e6965",
          6143 => x"642e0a00",
          6144 => x"46696c65",
          6145 => x"20616c72",
          6146 => x"65616479",
          6147 => x"20657869",
          6148 => x"7374732e",
          6149 => x"0a000000",
          6150 => x"46696c65",
          6151 => x"2068616e",
          6152 => x"646c6520",
          6153 => x"696e7661",
          6154 => x"6c69642e",
          6155 => x"0a000000",
          6156 => x"53442069",
          6157 => x"73207772",
          6158 => x"69746520",
          6159 => x"70726f74",
          6160 => x"65637465",
          6161 => x"642e0a00",
          6162 => x"44726976",
          6163 => x"65206e75",
          6164 => x"6d626572",
          6165 => x"20697320",
          6166 => x"696e7661",
          6167 => x"6c69642e",
          6168 => x"0a000000",
          6169 => x"4469736b",
          6170 => x"206e6f74",
          6171 => x"20656e61",
          6172 => x"626c6564",
          6173 => x"2e0a0000",
          6174 => x"4e6f2063",
          6175 => x"6f6d7061",
          6176 => x"7469626c",
          6177 => x"65206669",
          6178 => x"6c657379",
          6179 => x"7374656d",
          6180 => x"20666f75",
          6181 => x"6e64206f",
          6182 => x"6e206469",
          6183 => x"736b2e0a",
          6184 => x"00000000",
          6185 => x"466f726d",
          6186 => x"61742061",
          6187 => x"626f7274",
          6188 => x"65642e0a",
          6189 => x"00000000",
          6190 => x"54696d65",
          6191 => x"6f75742c",
          6192 => x"206f7065",
          6193 => x"72617469",
          6194 => x"6f6e2063",
          6195 => x"616e6365",
          6196 => x"6c6c6564",
          6197 => x"2e0a0000",
          6198 => x"46696c65",
          6199 => x"20697320",
          6200 => x"6c6f636b",
          6201 => x"65642e0a",
          6202 => x"00000000",
          6203 => x"496e7375",
          6204 => x"66666963",
          6205 => x"69656e74",
          6206 => x"206d656d",
          6207 => x"6f72792e",
          6208 => x"0a000000",
          6209 => x"546f6f20",
          6210 => x"6d616e79",
          6211 => x"206f7065",
          6212 => x"6e206669",
          6213 => x"6c65732e",
          6214 => x"0a000000",
          6215 => x"50617261",
          6216 => x"6d657465",
          6217 => x"72732069",
          6218 => x"6e636f72",
          6219 => x"72656374",
          6220 => x"2e0a0000",
          6221 => x"53756363",
          6222 => x"6573732e",
          6223 => x"0a000000",
          6224 => x"556e6b6e",
          6225 => x"6f776e20",
          6226 => x"6572726f",
          6227 => x"722e0a00",
          6228 => x"0a256c75",
          6229 => x"20627974",
          6230 => x"65732025",
          6231 => x"73206174",
          6232 => x"20256c75",
          6233 => x"20627974",
          6234 => x"65732f73",
          6235 => x"65632e0a",
          6236 => x"00000000",
          6237 => x"72656164",
          6238 => x"00000000",
          6239 => x"25303858",
          6240 => x"00000000",
          6241 => x"3a202000",
          6242 => x"25303458",
          6243 => x"00000000",
          6244 => x"20202020",
          6245 => x"20202020",
          6246 => x"00000000",
          6247 => x"25303258",
          6248 => x"00000000",
          6249 => x"20200000",
          6250 => x"207c0000",
          6251 => x"7c0d0a00",
          6252 => x"7a4f5300",
          6253 => x"0a2a2a20",
          6254 => x"25732028",
          6255 => x"00000000",
          6256 => x"31302f30",
          6257 => x"342f3230",
          6258 => x"32300000",
          6259 => x"76312e30",
          6260 => x"00000000",
          6261 => x"205a5055",
          6262 => x"2c207265",
          6263 => x"76202530",
          6264 => x"32782920",
          6265 => x"25732025",
          6266 => x"73202a2a",
          6267 => x"0a0a0000",
          6268 => x"5a505520",
          6269 => x"496e7465",
          6270 => x"72727570",
          6271 => x"74204861",
          6272 => x"6e646c65",
          6273 => x"720a0000",
          6274 => x"54696d65",
          6275 => x"7220696e",
          6276 => x"74657272",
          6277 => x"7570740a",
          6278 => x"00000000",
          6279 => x"50533220",
          6280 => x"696e7465",
          6281 => x"72727570",
          6282 => x"740a0000",
          6283 => x"494f4354",
          6284 => x"4c205244",
          6285 => x"20696e74",
          6286 => x"65727275",
          6287 => x"70740a00",
          6288 => x"494f4354",
          6289 => x"4c205752",
          6290 => x"20696e74",
          6291 => x"65727275",
          6292 => x"70740a00",
          6293 => x"55415254",
          6294 => x"30205258",
          6295 => x"20696e74",
          6296 => x"65727275",
          6297 => x"70740a00",
          6298 => x"55415254",
          6299 => x"30205458",
          6300 => x"20696e74",
          6301 => x"65727275",
          6302 => x"70740a00",
          6303 => x"55415254",
          6304 => x"31205258",
          6305 => x"20696e74",
          6306 => x"65727275",
          6307 => x"70740a00",
          6308 => x"55415254",
          6309 => x"31205458",
          6310 => x"20696e74",
          6311 => x"65727275",
          6312 => x"70740a00",
          6313 => x"53657474",
          6314 => x"696e6720",
          6315 => x"75702074",
          6316 => x"696d6572",
          6317 => x"2e2e2e0a",
          6318 => x"00000000",
          6319 => x"456e6162",
          6320 => x"6c696e67",
          6321 => x"2074696d",
          6322 => x"65722e2e",
          6323 => x"2e0a0000",
          6324 => x"6175746f",
          6325 => x"65786563",
          6326 => x"2e626174",
          6327 => x"00000000",
          6328 => x"303a0000",
          6329 => x"4661696c",
          6330 => x"65642074",
          6331 => x"6f20696e",
          6332 => x"69746961",
          6333 => x"6c697365",
          6334 => x"20736420",
          6335 => x"63617264",
          6336 => x"20302c20",
          6337 => x"706c6561",
          6338 => x"73652069",
          6339 => x"6e697420",
          6340 => x"6d616e75",
          6341 => x"616c6c79",
          6342 => x"2e0a0000",
          6343 => x"2a200000",
          6344 => x"436c6561",
          6345 => x"72696e67",
          6346 => x"2e2e2e2e",
          6347 => x"00000000",
          6348 => x"436f7079",
          6349 => x"696e672e",
          6350 => x"2e2e0000",
          6351 => x"436f6d70",
          6352 => x"6172696e",
          6353 => x"672e2e2e",
          6354 => x"00000000",
          6355 => x"2530386c",
          6356 => x"78282530",
          6357 => x"3878292d",
          6358 => x"3e253038",
          6359 => x"6c782825",
          6360 => x"30387829",
          6361 => x"0a000000",
          6362 => x"44756d70",
          6363 => x"204d656d",
          6364 => x"6f72790a",
          6365 => x"00000000",
          6366 => x"0a436f6d",
          6367 => x"706c6574",
          6368 => x"652e0a00",
          6369 => x"25303858",
          6370 => x"20253032",
          6371 => x"582d0000",
          6372 => x"3f3f3f0a",
          6373 => x"00000000",
          6374 => x"25303858",
          6375 => x"20253034",
          6376 => x"582d0000",
          6377 => x"25303858",
          6378 => x"20253038",
          6379 => x"582d0000",
          6380 => x"45786563",
          6381 => x"7574696e",
          6382 => x"6720636f",
          6383 => x"64652040",
          6384 => x"20253038",
          6385 => x"78202e2e",
          6386 => x"2e0a0000",
          6387 => x"43616c6c",
          6388 => x"696e6720",
          6389 => x"636f6465",
          6390 => x"20402025",
          6391 => x"30387820",
          6392 => x"2e2e2e0a",
          6393 => x"00000000",
          6394 => x"43616c6c",
          6395 => x"20726574",
          6396 => x"75726e65",
          6397 => x"6420636f",
          6398 => x"64652028",
          6399 => x"2564292e",
          6400 => x"0a000000",
          6401 => x"52657374",
          6402 => x"61727469",
          6403 => x"6e672061",
          6404 => x"70706c69",
          6405 => x"63617469",
          6406 => x"6f6e2e2e",
          6407 => x"2e0a0000",
          6408 => x"436f6c64",
          6409 => x"20726562",
          6410 => x"6f6f7469",
          6411 => x"6e672e2e",
          6412 => x"2e0a0000",
          6413 => x"5a505500",
          6414 => x"62696e00",
          6415 => x"25643a5c",
          6416 => x"25735c25",
          6417 => x"732e2573",
          6418 => x"00000000",
          6419 => x"25643a5c",
          6420 => x"25735c25",
          6421 => x"73000000",
          6422 => x"25643a5c",
          6423 => x"25730000",
          6424 => x"42616420",
          6425 => x"636f6d6d",
          6426 => x"616e642e",
          6427 => x"0a000000",
          6428 => x"52756e6e",
          6429 => x"696e672e",
          6430 => x"2e2e0a00",
          6431 => x"456e6162",
          6432 => x"6c696e67",
          6433 => x"20696e74",
          6434 => x"65727275",
          6435 => x"7074732e",
          6436 => x"2e2e0a00",
          6437 => x"00000000",
          6438 => x"00000000",
          6439 => x"00007fff",
          6440 => x"00000000",
          6441 => x"00007fff",
          6442 => x"00010000",
          6443 => x"00007fff",
          6444 => x"00010000",
          6445 => x"00810000",
          6446 => x"01000000",
          6447 => x"017fffff",
          6448 => x"00000000",
          6449 => x"00000000",
          6450 => x"00007800",
          6451 => x"00000000",
          6452 => x"05f5e100",
          6453 => x"05f5e100",
          6454 => x"05f5e100",
          6455 => x"00000000",
          6456 => x"01010101",
          6457 => x"01010101",
          6458 => x"01011001",
          6459 => x"01000000",
          6460 => x"00000000",
          6461 => x"01000000",
          6462 => x"00000000",
          6463 => x"00007ef0",
          6464 => x"01020100",
          6465 => x"00000000",
          6466 => x"00000000",
          6467 => x"00007ef8",
          6468 => x"01040100",
          6469 => x"00000000",
          6470 => x"00000000",
          6471 => x"00007f00",
          6472 => x"01140300",
          6473 => x"00000000",
          6474 => x"00000000",
          6475 => x"00007f08",
          6476 => x"012b0300",
          6477 => x"00000000",
          6478 => x"00000000",
          6479 => x"00007f10",
          6480 => x"01300300",
          6481 => x"00000000",
          6482 => x"00000000",
          6483 => x"00007f18",
          6484 => x"013c0400",
          6485 => x"00000000",
          6486 => x"00000000",
          6487 => x"00007f20",
          6488 => x"013d0400",
          6489 => x"00000000",
          6490 => x"00000000",
          6491 => x"00007f28",
          6492 => x"013f0400",
          6493 => x"00000000",
          6494 => x"00000000",
          6495 => x"00007f30",
          6496 => x"01400400",
          6497 => x"00000000",
          6498 => x"00000000",
          6499 => x"00007f38",
          6500 => x"01410400",
          6501 => x"00000000",
          6502 => x"00000000",
          6503 => x"00007f3c",
          6504 => x"01420400",
          6505 => x"00000000",
          6506 => x"00000000",
          6507 => x"00007f40",
          6508 => x"01430400",
          6509 => x"00000000",
          6510 => x"00000000",
          6511 => x"00007f44",
          6512 => x"01500500",
          6513 => x"00000000",
          6514 => x"00000000",
          6515 => x"00007f48",
          6516 => x"01510500",
          6517 => x"00000000",
          6518 => x"00000000",
          6519 => x"00007f4c",
          6520 => x"01540500",
          6521 => x"00000000",
          6522 => x"00000000",
          6523 => x"00007f50",
          6524 => x"01550500",
          6525 => x"00000000",
          6526 => x"00000000",
          6527 => x"00007f54",
          6528 => x"01790700",
          6529 => x"00000000",
          6530 => x"00000000",
          6531 => x"00007f5c",
          6532 => x"01780700",
          6533 => x"00000000",
          6534 => x"00000000",
          6535 => x"00007f60",
          6536 => x"01820800",
          6537 => x"00000000",
          6538 => x"00000000",
          6539 => x"00007f68",
          6540 => x"01830800",
          6541 => x"00000000",
          6542 => x"00000000",
          6543 => x"00007f70",
          6544 => x"01850800",
          6545 => x"00000000",
          6546 => x"00000000",
          6547 => x"00007f78",
          6548 => x"01870800",
          6549 => x"00000000",
          6550 => x"00000000",
          6551 => x"00007f80",
          6552 => x"018c0900",
          6553 => x"00000000",
          6554 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

