-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"b0",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"bd",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"ac",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"ab",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8f",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"90",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"91",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"92",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"f0",
           386 => x"ec",
           387 => x"f0",
           388 => x"80",
           389 => x"b8",
           390 => x"ee",
           391 => x"f0",
           392 => x"80",
           393 => x"b8",
           394 => x"f3",
           395 => x"f0",
           396 => x"80",
           397 => x"b8",
           398 => x"e0",
           399 => x"f0",
           400 => x"80",
           401 => x"b8",
           402 => x"a3",
           403 => x"f0",
           404 => x"80",
           405 => x"b8",
           406 => x"f6",
           407 => x"f0",
           408 => x"80",
           409 => x"b8",
           410 => x"86",
           411 => x"f0",
           412 => x"80",
           413 => x"b8",
           414 => x"82",
           415 => x"f0",
           416 => x"80",
           417 => x"b8",
           418 => x"88",
           419 => x"f0",
           420 => x"80",
           421 => x"b8",
           422 => x"a8",
           423 => x"f0",
           424 => x"80",
           425 => x"b8",
           426 => x"d1",
           427 => x"f0",
           428 => x"80",
           429 => x"b8",
           430 => x"8a",
           431 => x"f0",
           432 => x"80",
           433 => x"b8",
           434 => x"d4",
           435 => x"b8",
           436 => x"c0",
           437 => x"84",
           438 => x"80",
           439 => x"84",
           440 => x"80",
           441 => x"04",
           442 => x"0c",
           443 => x"2d",
           444 => x"08",
           445 => x"90",
           446 => x"f0",
           447 => x"c0",
           448 => x"f0",
           449 => x"80",
           450 => x"b8",
           451 => x"c9",
           452 => x"b8",
           453 => x"c0",
           454 => x"84",
           455 => x"82",
           456 => x"84",
           457 => x"80",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"90",
           463 => x"f0",
           464 => x"af",
           465 => x"f0",
           466 => x"80",
           467 => x"b8",
           468 => x"ed",
           469 => x"b8",
           470 => x"c0",
           471 => x"84",
           472 => x"82",
           473 => x"84",
           474 => x"80",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"90",
           480 => x"f0",
           481 => x"ad",
           482 => x"f0",
           483 => x"80",
           484 => x"b8",
           485 => x"f2",
           486 => x"b8",
           487 => x"c0",
           488 => x"84",
           489 => x"82",
           490 => x"84",
           491 => x"80",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"90",
           497 => x"f0",
           498 => x"d6",
           499 => x"f0",
           500 => x"80",
           501 => x"b8",
           502 => x"8a",
           503 => x"b8",
           504 => x"c0",
           505 => x"84",
           506 => x"82",
           507 => x"84",
           508 => x"80",
           509 => x"04",
           510 => x"0c",
           511 => x"2d",
           512 => x"08",
           513 => x"90",
           514 => x"f0",
           515 => x"f7",
           516 => x"f0",
           517 => x"80",
           518 => x"b8",
           519 => x"e5",
           520 => x"b8",
           521 => x"c0",
           522 => x"84",
           523 => x"82",
           524 => x"84",
           525 => x"80",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"90",
           531 => x"f0",
           532 => x"96",
           533 => x"f0",
           534 => x"80",
           535 => x"b8",
           536 => x"96",
           537 => x"b8",
           538 => x"c0",
           539 => x"84",
           540 => x"83",
           541 => x"84",
           542 => x"80",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"90",
           548 => x"f0",
           549 => x"ee",
           550 => x"f0",
           551 => x"80",
           552 => x"b8",
           553 => x"a4",
           554 => x"b8",
           555 => x"c0",
           556 => x"84",
           557 => x"83",
           558 => x"84",
           559 => x"80",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"90",
           565 => x"f0",
           566 => x"d2",
           567 => x"f0",
           568 => x"80",
           569 => x"b8",
           570 => x"f4",
           571 => x"b8",
           572 => x"c0",
           573 => x"84",
           574 => x"81",
           575 => x"84",
           576 => x"80",
           577 => x"04",
           578 => x"0c",
           579 => x"2d",
           580 => x"08",
           581 => x"90",
           582 => x"f0",
           583 => x"df",
           584 => x"f0",
           585 => x"80",
           586 => x"b8",
           587 => x"d7",
           588 => x"b8",
           589 => x"c0",
           590 => x"84",
           591 => x"b1",
           592 => x"b8",
           593 => x"c0",
           594 => x"84",
           595 => x"81",
           596 => x"84",
           597 => x"80",
           598 => x"04",
           599 => x"0c",
           600 => x"2d",
           601 => x"08",
           602 => x"90",
           603 => x"f0",
           604 => x"ac",
           605 => x"f0",
           606 => x"80",
           607 => x"b8",
           608 => x"d5",
           609 => x"b8",
           610 => x"c0",
           611 => x"3c",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"00",
           621 => x"ff",
           622 => x"06",
           623 => x"83",
           624 => x"10",
           625 => x"fc",
           626 => x"51",
           627 => x"80",
           628 => x"ff",
           629 => x"06",
           630 => x"52",
           631 => x"0a",
           632 => x"38",
           633 => x"51",
           634 => x"e4",
           635 => x"d0",
           636 => x"80",
           637 => x"05",
           638 => x"0b",
           639 => x"04",
           640 => x"80",
           641 => x"00",
           642 => x"87",
           643 => x"84",
           644 => x"56",
           645 => x"84",
           646 => x"51",
           647 => x"86",
           648 => x"fa",
           649 => x"7a",
           650 => x"33",
           651 => x"06",
           652 => x"07",
           653 => x"57",
           654 => x"72",
           655 => x"06",
           656 => x"ff",
           657 => x"8a",
           658 => x"70",
           659 => x"2a",
           660 => x"56",
           661 => x"25",
           662 => x"80",
           663 => x"75",
           664 => x"3f",
           665 => x"08",
           666 => x"e4",
           667 => x"ae",
           668 => x"e4",
           669 => x"81",
           670 => x"ff",
           671 => x"32",
           672 => x"72",
           673 => x"51",
           674 => x"73",
           675 => x"38",
           676 => x"76",
           677 => x"b8",
           678 => x"3d",
           679 => x"0b",
           680 => x"0c",
           681 => x"04",
           682 => x"7d",
           683 => x"84",
           684 => x"34",
           685 => x"0a",
           686 => x"88",
           687 => x"52",
           688 => x"05",
           689 => x"73",
           690 => x"74",
           691 => x"0d",
           692 => x"0d",
           693 => x"05",
           694 => x"75",
           695 => x"85",
           696 => x"f1",
           697 => x"63",
           698 => x"5d",
           699 => x"1f",
           700 => x"33",
           701 => x"81",
           702 => x"55",
           703 => x"54",
           704 => x"09",
           705 => x"d2",
           706 => x"57",
           707 => x"80",
           708 => x"1c",
           709 => x"54",
           710 => x"2e",
           711 => x"d0",
           712 => x"89",
           713 => x"38",
           714 => x"70",
           715 => x"25",
           716 => x"78",
           717 => x"80",
           718 => x"7a",
           719 => x"81",
           720 => x"40",
           721 => x"2e",
           722 => x"82",
           723 => x"7b",
           724 => x"ff",
           725 => x"1d",
           726 => x"84",
           727 => x"91",
           728 => x"7a",
           729 => x"78",
           730 => x"79",
           731 => x"98",
           732 => x"2c",
           733 => x"80",
           734 => x"0a",
           735 => x"2c",
           736 => x"56",
           737 => x"24",
           738 => x"73",
           739 => x"72",
           740 => x"78",
           741 => x"58",
           742 => x"38",
           743 => x"76",
           744 => x"81",
           745 => x"81",
           746 => x"5a",
           747 => x"33",
           748 => x"fe",
           749 => x"9e",
           750 => x"76",
           751 => x"3f",
           752 => x"76",
           753 => x"ff",
           754 => x"83",
           755 => x"06",
           756 => x"8a",
           757 => x"74",
           758 => x"7e",
           759 => x"17",
           760 => x"d8",
           761 => x"72",
           762 => x"c9",
           763 => x"73",
           764 => x"e0",
           765 => x"80",
           766 => x"eb",
           767 => x"76",
           768 => x"3f",
           769 => x"58",
           770 => x"86",
           771 => x"39",
           772 => x"fe",
           773 => x"5a",
           774 => x"05",
           775 => x"83",
           776 => x"5e",
           777 => x"84",
           778 => x"79",
           779 => x"93",
           780 => x"b8",
           781 => x"ff",
           782 => x"e4",
           783 => x"05",
           784 => x"89",
           785 => x"84",
           786 => x"b0",
           787 => x"7e",
           788 => x"40",
           789 => x"75",
           790 => x"3f",
           791 => x"08",
           792 => x"e4",
           793 => x"7d",
           794 => x"31",
           795 => x"b2",
           796 => x"7e",
           797 => x"38",
           798 => x"80",
           799 => x"80",
           800 => x"2c",
           801 => x"86",
           802 => x"06",
           803 => x"80",
           804 => x"77",
           805 => x"29",
           806 => x"05",
           807 => x"2e",
           808 => x"84",
           809 => x"fc",
           810 => x"53",
           811 => x"58",
           812 => x"70",
           813 => x"55",
           814 => x"9e",
           815 => x"2c",
           816 => x"06",
           817 => x"73",
           818 => x"38",
           819 => x"f7",
           820 => x"2a",
           821 => x"41",
           822 => x"81",
           823 => x"80",
           824 => x"38",
           825 => x"90",
           826 => x"2c",
           827 => x"06",
           828 => x"73",
           829 => x"96",
           830 => x"2a",
           831 => x"73",
           832 => x"7a",
           833 => x"06",
           834 => x"98",
           835 => x"2a",
           836 => x"73",
           837 => x"7e",
           838 => x"73",
           839 => x"7a",
           840 => x"06",
           841 => x"2e",
           842 => x"78",
           843 => x"29",
           844 => x"05",
           845 => x"5a",
           846 => x"74",
           847 => x"7c",
           848 => x"88",
           849 => x"78",
           850 => x"29",
           851 => x"05",
           852 => x"5a",
           853 => x"80",
           854 => x"74",
           855 => x"72",
           856 => x"38",
           857 => x"80",
           858 => x"ff",
           859 => x"98",
           860 => x"55",
           861 => x"9d",
           862 => x"b0",
           863 => x"3f",
           864 => x"80",
           865 => x"ff",
           866 => x"98",
           867 => x"55",
           868 => x"e5",
           869 => x"2a",
           870 => x"5c",
           871 => x"2e",
           872 => x"76",
           873 => x"84",
           874 => x"80",
           875 => x"ca",
           876 => x"d3",
           877 => x"38",
           878 => x"f4",
           879 => x"7c",
           880 => x"70",
           881 => x"87",
           882 => x"84",
           883 => x"09",
           884 => x"38",
           885 => x"5b",
           886 => x"fc",
           887 => x"78",
           888 => x"29",
           889 => x"05",
           890 => x"5a",
           891 => x"75",
           892 => x"38",
           893 => x"51",
           894 => x"e2",
           895 => x"07",
           896 => x"07",
           897 => x"5b",
           898 => x"38",
           899 => x"7a",
           900 => x"5b",
           901 => x"90",
           902 => x"05",
           903 => x"83",
           904 => x"5f",
           905 => x"5a",
           906 => x"7f",
           907 => x"77",
           908 => x"06",
           909 => x"70",
           910 => x"07",
           911 => x"80",
           912 => x"80",
           913 => x"2c",
           914 => x"56",
           915 => x"7a",
           916 => x"81",
           917 => x"7a",
           918 => x"77",
           919 => x"80",
           920 => x"80",
           921 => x"2c",
           922 => x"80",
           923 => x"b3",
           924 => x"a0",
           925 => x"3f",
           926 => x"1a",
           927 => x"ff",
           928 => x"79",
           929 => x"2e",
           930 => x"7c",
           931 => x"81",
           932 => x"51",
           933 => x"e2",
           934 => x"70",
           935 => x"06",
           936 => x"83",
           937 => x"fe",
           938 => x"52",
           939 => x"05",
           940 => x"85",
           941 => x"39",
           942 => x"06",
           943 => x"07",
           944 => x"80",
           945 => x"80",
           946 => x"2c",
           947 => x"80",
           948 => x"2a",
           949 => x"5d",
           950 => x"fd",
           951 => x"fb",
           952 => x"84",
           953 => x"70",
           954 => x"56",
           955 => x"82",
           956 => x"83",
           957 => x"5b",
           958 => x"5e",
           959 => x"7a",
           960 => x"33",
           961 => x"f8",
           962 => x"ca",
           963 => x"07",
           964 => x"33",
           965 => x"f7",
           966 => x"ba",
           967 => x"84",
           968 => x"77",
           969 => x"58",
           970 => x"82",
           971 => x"51",
           972 => x"84",
           973 => x"83",
           974 => x"78",
           975 => x"2b",
           976 => x"90",
           977 => x"87",
           978 => x"c0",
           979 => x"58",
           980 => x"be",
           981 => x"39",
           982 => x"05",
           983 => x"81",
           984 => x"41",
           985 => x"cf",
           986 => x"87",
           987 => x"b8",
           988 => x"ff",
           989 => x"71",
           990 => x"54",
           991 => x"7a",
           992 => x"7c",
           993 => x"76",
           994 => x"f7",
           995 => x"78",
           996 => x"29",
           997 => x"05",
           998 => x"5a",
           999 => x"74",
          1000 => x"38",
          1001 => x"51",
          1002 => x"e2",
          1003 => x"b0",
          1004 => x"3f",
          1005 => x"09",
          1006 => x"e3",
          1007 => x"76",
          1008 => x"3f",
          1009 => x"81",
          1010 => x"80",
          1011 => x"38",
          1012 => x"75",
          1013 => x"71",
          1014 => x"70",
          1015 => x"83",
          1016 => x"5a",
          1017 => x"fa",
          1018 => x"a2",
          1019 => x"ad",
          1020 => x"3f",
          1021 => x"54",
          1022 => x"fa",
          1023 => x"ad",
          1024 => x"75",
          1025 => x"82",
          1026 => x"81",
          1027 => x"80",
          1028 => x"38",
          1029 => x"78",
          1030 => x"2b",
          1031 => x"5a",
          1032 => x"39",
          1033 => x"51",
          1034 => x"c8",
          1035 => x"a0",
          1036 => x"3f",
          1037 => x"78",
          1038 => x"88",
          1039 => x"b8",
          1040 => x"ff",
          1041 => x"71",
          1042 => x"54",
          1043 => x"39",
          1044 => x"7e",
          1045 => x"ff",
          1046 => x"57",
          1047 => x"39",
          1048 => x"84",
          1049 => x"53",
          1050 => x"51",
          1051 => x"84",
          1052 => x"fa",
          1053 => x"55",
          1054 => x"d4",
          1055 => x"11",
          1056 => x"2a",
          1057 => x"81",
          1058 => x"58",
          1059 => x"56",
          1060 => x"09",
          1061 => x"d5",
          1062 => x"81",
          1063 => x"53",
          1064 => x"b0",
          1065 => x"c8",
          1066 => x"51",
          1067 => x"53",
          1068 => x"b8",
          1069 => x"2e",
          1070 => x"57",
          1071 => x"05",
          1072 => x"72",
          1073 => x"38",
          1074 => x"08",
          1075 => x"84",
          1076 => x"54",
          1077 => x"08",
          1078 => x"90",
          1079 => x"74",
          1080 => x"e4",
          1081 => x"83",
          1082 => x"76",
          1083 => x"b8",
          1084 => x"3d",
          1085 => x"3d",
          1086 => x"56",
          1087 => x"85",
          1088 => x"81",
          1089 => x"70",
          1090 => x"55",
          1091 => x"56",
          1092 => x"09",
          1093 => x"38",
          1094 => x"05",
          1095 => x"72",
          1096 => x"81",
          1097 => x"76",
          1098 => x"b8",
          1099 => x"3d",
          1100 => x"70",
          1101 => x"33",
          1102 => x"2e",
          1103 => x"52",
          1104 => x"15",
          1105 => x"2d",
          1106 => x"08",
          1107 => x"38",
          1108 => x"81",
          1109 => x"54",
          1110 => x"38",
          1111 => x"3d",
          1112 => x"c8",
          1113 => x"51",
          1114 => x"3d",
          1115 => x"3d",
          1116 => x"85",
          1117 => x"81",
          1118 => x"81",
          1119 => x"56",
          1120 => x"72",
          1121 => x"82",
          1122 => x"54",
          1123 => x"ac",
          1124 => x"08",
          1125 => x"16",
          1126 => x"38",
          1127 => x"76",
          1128 => x"08",
          1129 => x"0c",
          1130 => x"53",
          1131 => x"16",
          1132 => x"75",
          1133 => x"0c",
          1134 => x"04",
          1135 => x"81",
          1136 => x"90",
          1137 => x"73",
          1138 => x"84",
          1139 => x"e3",
          1140 => x"08",
          1141 => x"16",
          1142 => x"d7",
          1143 => x"0d",
          1144 => x"33",
          1145 => x"06",
          1146 => x"81",
          1147 => x"56",
          1148 => x"71",
          1149 => x"86",
          1150 => x"52",
          1151 => x"72",
          1152 => x"06",
          1153 => x"2e",
          1154 => x"75",
          1155 => x"53",
          1156 => x"2e",
          1157 => x"81",
          1158 => x"8c",
          1159 => x"05",
          1160 => x"71",
          1161 => x"54",
          1162 => x"e4",
          1163 => x"0d",
          1164 => x"bf",
          1165 => x"85",
          1166 => x"16",
          1167 => x"8c",
          1168 => x"16",
          1169 => x"e4",
          1170 => x"0d",
          1171 => x"94",
          1172 => x"74",
          1173 => x"e4",
          1174 => x"b8",
          1175 => x"25",
          1176 => x"85",
          1177 => x"90",
          1178 => x"84",
          1179 => x"ff",
          1180 => x"71",
          1181 => x"72",
          1182 => x"ff",
          1183 => x"b8",
          1184 => x"3d",
          1185 => x"a0",
          1186 => x"85",
          1187 => x"54",
          1188 => x"3d",
          1189 => x"71",
          1190 => x"71",
          1191 => x"53",
          1192 => x"f7",
          1193 => x"52",
          1194 => x"05",
          1195 => x"70",
          1196 => x"05",
          1197 => x"f0",
          1198 => x"b8",
          1199 => x"3d",
          1200 => x"3d",
          1201 => x"71",
          1202 => x"52",
          1203 => x"2e",
          1204 => x"72",
          1205 => x"70",
          1206 => x"38",
          1207 => x"05",
          1208 => x"70",
          1209 => x"34",
          1210 => x"70",
          1211 => x"84",
          1212 => x"86",
          1213 => x"70",
          1214 => x"75",
          1215 => x"70",
          1216 => x"53",
          1217 => x"13",
          1218 => x"33",
          1219 => x"11",
          1220 => x"2e",
          1221 => x"13",
          1222 => x"53",
          1223 => x"34",
          1224 => x"70",
          1225 => x"39",
          1226 => x"74",
          1227 => x"71",
          1228 => x"53",
          1229 => x"f7",
          1230 => x"70",
          1231 => x"b8",
          1232 => x"84",
          1233 => x"fd",
          1234 => x"77",
          1235 => x"54",
          1236 => x"05",
          1237 => x"70",
          1238 => x"05",
          1239 => x"f0",
          1240 => x"b8",
          1241 => x"3d",
          1242 => x"3d",
          1243 => x"71",
          1244 => x"52",
          1245 => x"2e",
          1246 => x"70",
          1247 => x"33",
          1248 => x"05",
          1249 => x"11",
          1250 => x"38",
          1251 => x"e4",
          1252 => x"0d",
          1253 => x"0d",
          1254 => x"55",
          1255 => x"80",
          1256 => x"73",
          1257 => x"81",
          1258 => x"52",
          1259 => x"2e",
          1260 => x"9a",
          1261 => x"54",
          1262 => x"b7",
          1263 => x"53",
          1264 => x"80",
          1265 => x"b8",
          1266 => x"3d",
          1267 => x"80",
          1268 => x"73",
          1269 => x"51",
          1270 => x"e9",
          1271 => x"33",
          1272 => x"71",
          1273 => x"38",
          1274 => x"84",
          1275 => x"86",
          1276 => x"71",
          1277 => x"0c",
          1278 => x"04",
          1279 => x"77",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"08",
          1284 => x"55",
          1285 => x"3f",
          1286 => x"08",
          1287 => x"e4",
          1288 => x"9b",
          1289 => x"e4",
          1290 => x"80",
          1291 => x"53",
          1292 => x"b8",
          1293 => x"fe",
          1294 => x"b8",
          1295 => x"73",
          1296 => x"0c",
          1297 => x"04",
          1298 => x"75",
          1299 => x"54",
          1300 => x"71",
          1301 => x"38",
          1302 => x"05",
          1303 => x"70",
          1304 => x"38",
          1305 => x"71",
          1306 => x"81",
          1307 => x"ff",
          1308 => x"31",
          1309 => x"84",
          1310 => x"85",
          1311 => x"fd",
          1312 => x"77",
          1313 => x"53",
          1314 => x"80",
          1315 => x"72",
          1316 => x"05",
          1317 => x"11",
          1318 => x"38",
          1319 => x"e4",
          1320 => x"0d",
          1321 => x"0d",
          1322 => x"54",
          1323 => x"80",
          1324 => x"76",
          1325 => x"3f",
          1326 => x"08",
          1327 => x"53",
          1328 => x"8d",
          1329 => x"80",
          1330 => x"84",
          1331 => x"31",
          1332 => x"72",
          1333 => x"cb",
          1334 => x"72",
          1335 => x"c3",
          1336 => x"74",
          1337 => x"72",
          1338 => x"2b",
          1339 => x"55",
          1340 => x"76",
          1341 => x"72",
          1342 => x"2a",
          1343 => x"77",
          1344 => x"31",
          1345 => x"2c",
          1346 => x"7b",
          1347 => x"71",
          1348 => x"5c",
          1349 => x"55",
          1350 => x"74",
          1351 => x"10",
          1352 => x"71",
          1353 => x"0c",
          1354 => x"04",
          1355 => x"76",
          1356 => x"80",
          1357 => x"70",
          1358 => x"25",
          1359 => x"90",
          1360 => x"71",
          1361 => x"fe",
          1362 => x"30",
          1363 => x"83",
          1364 => x"31",
          1365 => x"70",
          1366 => x"70",
          1367 => x"25",
          1368 => x"71",
          1369 => x"2a",
          1370 => x"1b",
          1371 => x"06",
          1372 => x"80",
          1373 => x"71",
          1374 => x"2a",
          1375 => x"81",
          1376 => x"06",
          1377 => x"74",
          1378 => x"19",
          1379 => x"e4",
          1380 => x"54",
          1381 => x"56",
          1382 => x"55",
          1383 => x"56",
          1384 => x"58",
          1385 => x"86",
          1386 => x"fd",
          1387 => x"77",
          1388 => x"53",
          1389 => x"94",
          1390 => x"e4",
          1391 => x"74",
          1392 => x"b8",
          1393 => x"85",
          1394 => x"fa",
          1395 => x"7a",
          1396 => x"53",
          1397 => x"8b",
          1398 => x"fe",
          1399 => x"b8",
          1400 => x"e0",
          1401 => x"80",
          1402 => x"73",
          1403 => x"3f",
          1404 => x"e4",
          1405 => x"73",
          1406 => x"26",
          1407 => x"80",
          1408 => x"2e",
          1409 => x"12",
          1410 => x"a0",
          1411 => x"71",
          1412 => x"54",
          1413 => x"74",
          1414 => x"38",
          1415 => x"9f",
          1416 => x"10",
          1417 => x"72",
          1418 => x"9f",
          1419 => x"06",
          1420 => x"75",
          1421 => x"1c",
          1422 => x"52",
          1423 => x"53",
          1424 => x"72",
          1425 => x"0c",
          1426 => x"04",
          1427 => x"78",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"9f",
          1431 => x"73",
          1432 => x"74",
          1433 => x"75",
          1434 => x"56",
          1435 => x"fc",
          1436 => x"b8",
          1437 => x"32",
          1438 => x"b8",
          1439 => x"3d",
          1440 => x"3d",
          1441 => x"5b",
          1442 => x"7b",
          1443 => x"70",
          1444 => x"59",
          1445 => x"09",
          1446 => x"38",
          1447 => x"78",
          1448 => x"55",
          1449 => x"2e",
          1450 => x"ad",
          1451 => x"38",
          1452 => x"81",
          1453 => x"14",
          1454 => x"77",
          1455 => x"db",
          1456 => x"80",
          1457 => x"27",
          1458 => x"80",
          1459 => x"89",
          1460 => x"70",
          1461 => x"55",
          1462 => x"70",
          1463 => x"51",
          1464 => x"27",
          1465 => x"13",
          1466 => x"06",
          1467 => x"73",
          1468 => x"38",
          1469 => x"81",
          1470 => x"76",
          1471 => x"16",
          1472 => x"70",
          1473 => x"56",
          1474 => x"ff",
          1475 => x"80",
          1476 => x"75",
          1477 => x"7a",
          1478 => x"75",
          1479 => x"0c",
          1480 => x"04",
          1481 => x"70",
          1482 => x"33",
          1483 => x"73",
          1484 => x"81",
          1485 => x"38",
          1486 => x"78",
          1487 => x"55",
          1488 => x"e2",
          1489 => x"90",
          1490 => x"f8",
          1491 => x"81",
          1492 => x"27",
          1493 => x"14",
          1494 => x"88",
          1495 => x"27",
          1496 => x"75",
          1497 => x"0c",
          1498 => x"04",
          1499 => x"15",
          1500 => x"70",
          1501 => x"80",
          1502 => x"39",
          1503 => x"b8",
          1504 => x"3d",
          1505 => x"3d",
          1506 => x"5b",
          1507 => x"7b",
          1508 => x"70",
          1509 => x"59",
          1510 => x"09",
          1511 => x"38",
          1512 => x"78",
          1513 => x"55",
          1514 => x"2e",
          1515 => x"ad",
          1516 => x"38",
          1517 => x"81",
          1518 => x"14",
          1519 => x"77",
          1520 => x"db",
          1521 => x"80",
          1522 => x"27",
          1523 => x"80",
          1524 => x"89",
          1525 => x"70",
          1526 => x"55",
          1527 => x"70",
          1528 => x"51",
          1529 => x"27",
          1530 => x"13",
          1531 => x"06",
          1532 => x"73",
          1533 => x"38",
          1534 => x"81",
          1535 => x"76",
          1536 => x"16",
          1537 => x"70",
          1538 => x"56",
          1539 => x"ff",
          1540 => x"80",
          1541 => x"75",
          1542 => x"7a",
          1543 => x"75",
          1544 => x"0c",
          1545 => x"04",
          1546 => x"70",
          1547 => x"33",
          1548 => x"73",
          1549 => x"81",
          1550 => x"38",
          1551 => x"78",
          1552 => x"55",
          1553 => x"e2",
          1554 => x"90",
          1555 => x"f8",
          1556 => x"81",
          1557 => x"27",
          1558 => x"14",
          1559 => x"88",
          1560 => x"27",
          1561 => x"75",
          1562 => x"0c",
          1563 => x"04",
          1564 => x"15",
          1565 => x"70",
          1566 => x"80",
          1567 => x"39",
          1568 => x"b8",
          1569 => x"3d",
          1570 => x"d6",
          1571 => x"b8",
          1572 => x"ff",
          1573 => x"e4",
          1574 => x"3d",
          1575 => x"71",
          1576 => x"38",
          1577 => x"83",
          1578 => x"52",
          1579 => x"83",
          1580 => x"ef",
          1581 => x"3d",
          1582 => x"ce",
          1583 => x"b3",
          1584 => x"0d",
          1585 => x"b4",
          1586 => x"3f",
          1587 => x"04",
          1588 => x"51",
          1589 => x"83",
          1590 => x"83",
          1591 => x"ef",
          1592 => x"3d",
          1593 => x"ce",
          1594 => x"87",
          1595 => x"0d",
          1596 => x"94",
          1597 => x"3f",
          1598 => x"04",
          1599 => x"51",
          1600 => x"83",
          1601 => x"83",
          1602 => x"ee",
          1603 => x"3d",
          1604 => x"cf",
          1605 => x"db",
          1606 => x"0d",
          1607 => x"fc",
          1608 => x"3f",
          1609 => x"04",
          1610 => x"51",
          1611 => x"83",
          1612 => x"83",
          1613 => x"ee",
          1614 => x"3d",
          1615 => x"d0",
          1616 => x"af",
          1617 => x"0d",
          1618 => x"d4",
          1619 => x"3f",
          1620 => x"04",
          1621 => x"51",
          1622 => x"83",
          1623 => x"83",
          1624 => x"ee",
          1625 => x"3d",
          1626 => x"d1",
          1627 => x"83",
          1628 => x"0d",
          1629 => x"98",
          1630 => x"3f",
          1631 => x"04",
          1632 => x"51",
          1633 => x"83",
          1634 => x"83",
          1635 => x"ed",
          1636 => x"3d",
          1637 => x"3d",
          1638 => x"84",
          1639 => x"05",
          1640 => x"80",
          1641 => x"70",
          1642 => x"25",
          1643 => x"59",
          1644 => x"87",
          1645 => x"38",
          1646 => x"77",
          1647 => x"ff",
          1648 => x"93",
          1649 => x"e2",
          1650 => x"77",
          1651 => x"70",
          1652 => x"95",
          1653 => x"b8",
          1654 => x"84",
          1655 => x"80",
          1656 => x"38",
          1657 => x"af",
          1658 => x"30",
          1659 => x"80",
          1660 => x"70",
          1661 => x"06",
          1662 => x"58",
          1663 => x"aa",
          1664 => x"98",
          1665 => x"74",
          1666 => x"80",
          1667 => x"52",
          1668 => x"29",
          1669 => x"3f",
          1670 => x"08",
          1671 => x"e4",
          1672 => x"83",
          1673 => x"df",
          1674 => x"84",
          1675 => x"96",
          1676 => x"84",
          1677 => x"87",
          1678 => x"0c",
          1679 => x"08",
          1680 => x"d4",
          1681 => x"80",
          1682 => x"77",
          1683 => x"bd",
          1684 => x"e4",
          1685 => x"b8",
          1686 => x"88",
          1687 => x"74",
          1688 => x"80",
          1689 => x"75",
          1690 => x"d5",
          1691 => x"52",
          1692 => x"b1",
          1693 => x"e4",
          1694 => x"51",
          1695 => x"84",
          1696 => x"54",
          1697 => x"53",
          1698 => x"d1",
          1699 => x"f8",
          1700 => x"39",
          1701 => x"7c",
          1702 => x"b7",
          1703 => x"59",
          1704 => x"53",
          1705 => x"51",
          1706 => x"84",
          1707 => x"8b",
          1708 => x"2e",
          1709 => x"81",
          1710 => x"77",
          1711 => x"0c",
          1712 => x"04",
          1713 => x"d4",
          1714 => x"55",
          1715 => x"b8",
          1716 => x"52",
          1717 => x"2d",
          1718 => x"08",
          1719 => x"0c",
          1720 => x"04",
          1721 => x"7f",
          1722 => x"8c",
          1723 => x"05",
          1724 => x"15",
          1725 => x"5c",
          1726 => x"5e",
          1727 => x"83",
          1728 => x"52",
          1729 => x"51",
          1730 => x"83",
          1731 => x"dd",
          1732 => x"54",
          1733 => x"b2",
          1734 => x"2e",
          1735 => x"7c",
          1736 => x"a8",
          1737 => x"53",
          1738 => x"81",
          1739 => x"33",
          1740 => x"f8",
          1741 => x"3f",
          1742 => x"d4",
          1743 => x"54",
          1744 => x"aa",
          1745 => x"26",
          1746 => x"d2",
          1747 => x"b8",
          1748 => x"75",
          1749 => x"c0",
          1750 => x"70",
          1751 => x"80",
          1752 => x"27",
          1753 => x"55",
          1754 => x"74",
          1755 => x"81",
          1756 => x"06",
          1757 => x"06",
          1758 => x"80",
          1759 => x"80",
          1760 => x"81",
          1761 => x"d4",
          1762 => x"a0",
          1763 => x"3f",
          1764 => x"78",
          1765 => x"38",
          1766 => x"51",
          1767 => x"78",
          1768 => x"5c",
          1769 => x"9d",
          1770 => x"b8",
          1771 => x"2b",
          1772 => x"58",
          1773 => x"2e",
          1774 => x"76",
          1775 => x"c3",
          1776 => x"57",
          1777 => x"fe",
          1778 => x"0b",
          1779 => x"0c",
          1780 => x"04",
          1781 => x"51",
          1782 => x"81",
          1783 => x"c8",
          1784 => x"a0",
          1785 => x"3f",
          1786 => x"fe",
          1787 => x"da",
          1788 => x"98",
          1789 => x"3f",
          1790 => x"d4",
          1791 => x"54",
          1792 => x"ea",
          1793 => x"27",
          1794 => x"73",
          1795 => x"7a",
          1796 => x"72",
          1797 => x"d2",
          1798 => x"ec",
          1799 => x"84",
          1800 => x"53",
          1801 => x"ea",
          1802 => x"74",
          1803 => x"fe",
          1804 => x"d2",
          1805 => x"d0",
          1806 => x"84",
          1807 => x"53",
          1808 => x"ea",
          1809 => x"79",
          1810 => x"38",
          1811 => x"72",
          1812 => x"38",
          1813 => x"83",
          1814 => x"db",
          1815 => x"14",
          1816 => x"08",
          1817 => x"51",
          1818 => x"78",
          1819 => x"38",
          1820 => x"84",
          1821 => x"52",
          1822 => x"f2",
          1823 => x"56",
          1824 => x"80",
          1825 => x"84",
          1826 => x"81",
          1827 => x"88",
          1828 => x"2e",
          1829 => x"a0",
          1830 => x"d0",
          1831 => x"06",
          1832 => x"90",
          1833 => x"39",
          1834 => x"a5",
          1835 => x"e4",
          1836 => x"70",
          1837 => x"a0",
          1838 => x"72",
          1839 => x"30",
          1840 => x"73",
          1841 => x"51",
          1842 => x"57",
          1843 => x"80",
          1844 => x"38",
          1845 => x"f9",
          1846 => x"e4",
          1847 => x"70",
          1848 => x"a0",
          1849 => x"72",
          1850 => x"30",
          1851 => x"73",
          1852 => x"51",
          1853 => x"57",
          1854 => x"73",
          1855 => x"38",
          1856 => x"80",
          1857 => x"e4",
          1858 => x"0d",
          1859 => x"0d",
          1860 => x"80",
          1861 => x"c7",
          1862 => x"9c",
          1863 => x"d2",
          1864 => x"fe",
          1865 => x"9c",
          1866 => x"81",
          1867 => x"06",
          1868 => x"82",
          1869 => x"82",
          1870 => x"06",
          1871 => x"82",
          1872 => x"83",
          1873 => x"06",
          1874 => x"81",
          1875 => x"84",
          1876 => x"06",
          1877 => x"81",
          1878 => x"85",
          1879 => x"06",
          1880 => x"80",
          1881 => x"86",
          1882 => x"06",
          1883 => x"80",
          1884 => x"87",
          1885 => x"06",
          1886 => x"a9",
          1887 => x"2a",
          1888 => x"72",
          1889 => x"df",
          1890 => x"0d",
          1891 => x"9b",
          1892 => x"d2",
          1893 => x"8a",
          1894 => x"9b",
          1895 => x"c7",
          1896 => x"0d",
          1897 => x"9b",
          1898 => x"d3",
          1899 => x"f2",
          1900 => x"9b",
          1901 => x"88",
          1902 => x"53",
          1903 => x"c6",
          1904 => x"81",
          1905 => x"3f",
          1906 => x"51",
          1907 => x"80",
          1908 => x"3f",
          1909 => x"70",
          1910 => x"52",
          1911 => x"ff",
          1912 => x"39",
          1913 => x"a2",
          1914 => x"b0",
          1915 => x"3f",
          1916 => x"96",
          1917 => x"2a",
          1918 => x"51",
          1919 => x"2e",
          1920 => x"ff",
          1921 => x"51",
          1922 => x"83",
          1923 => x"9b",
          1924 => x"51",
          1925 => x"72",
          1926 => x"81",
          1927 => x"71",
          1928 => x"c2",
          1929 => x"39",
          1930 => x"de",
          1931 => x"d8",
          1932 => x"3f",
          1933 => x"d2",
          1934 => x"2a",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"ff",
          1938 => x"51",
          1939 => x"83",
          1940 => x"9a",
          1941 => x"51",
          1942 => x"72",
          1943 => x"81",
          1944 => x"71",
          1945 => x"e6",
          1946 => x"39",
          1947 => x"9a",
          1948 => x"fc",
          1949 => x"3f",
          1950 => x"8e",
          1951 => x"2a",
          1952 => x"51",
          1953 => x"2e",
          1954 => x"ff",
          1955 => x"3d",
          1956 => x"41",
          1957 => x"84",
          1958 => x"42",
          1959 => x"51",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"9b",
          1963 => x"78",
          1964 => x"b1",
          1965 => x"d0",
          1966 => x"3f",
          1967 => x"83",
          1968 => x"d6",
          1969 => x"48",
          1970 => x"80",
          1971 => x"eb",
          1972 => x"0b",
          1973 => x"33",
          1974 => x"06",
          1975 => x"80",
          1976 => x"38",
          1977 => x"83",
          1978 => x"81",
          1979 => x"7d",
          1980 => x"c1",
          1981 => x"5a",
          1982 => x"2e",
          1983 => x"79",
          1984 => x"a0",
          1985 => x"06",
          1986 => x"1a",
          1987 => x"5a",
          1988 => x"f6",
          1989 => x"7b",
          1990 => x"38",
          1991 => x"83",
          1992 => x"70",
          1993 => x"e7",
          1994 => x"b8",
          1995 => x"b8",
          1996 => x"7a",
          1997 => x"52",
          1998 => x"3f",
          1999 => x"08",
          2000 => x"1b",
          2001 => x"81",
          2002 => x"38",
          2003 => x"81",
          2004 => x"5b",
          2005 => x"c4",
          2006 => x"33",
          2007 => x"2e",
          2008 => x"80",
          2009 => x"51",
          2010 => x"84",
          2011 => x"5e",
          2012 => x"08",
          2013 => x"c9",
          2014 => x"e4",
          2015 => x"3d",
          2016 => x"51",
          2017 => x"84",
          2018 => x"60",
          2019 => x"5c",
          2020 => x"81",
          2021 => x"b8",
          2022 => x"e7",
          2023 => x"b8",
          2024 => x"26",
          2025 => x"81",
          2026 => x"5e",
          2027 => x"2e",
          2028 => x"7a",
          2029 => x"e2",
          2030 => x"2e",
          2031 => x"7b",
          2032 => x"83",
          2033 => x"7c",
          2034 => x"3f",
          2035 => x"58",
          2036 => x"57",
          2037 => x"55",
          2038 => x"80",
          2039 => x"80",
          2040 => x"51",
          2041 => x"84",
          2042 => x"84",
          2043 => x"09",
          2044 => x"72",
          2045 => x"51",
          2046 => x"80",
          2047 => x"26",
          2048 => x"5a",
          2049 => x"59",
          2050 => x"8d",
          2051 => x"70",
          2052 => x"5c",
          2053 => x"95",
          2054 => x"32",
          2055 => x"07",
          2056 => x"ee",
          2057 => x"2e",
          2058 => x"7d",
          2059 => x"d0",
          2060 => x"88",
          2061 => x"3f",
          2062 => x"f8",
          2063 => x"7e",
          2064 => x"3f",
          2065 => x"ed",
          2066 => x"81",
          2067 => x"59",
          2068 => x"38",
          2069 => x"d4",
          2070 => x"cf",
          2071 => x"88",
          2072 => x"b8",
          2073 => x"c5",
          2074 => x"0b",
          2075 => x"d8",
          2076 => x"f4",
          2077 => x"52",
          2078 => x"f6",
          2079 => x"b8",
          2080 => x"2e",
          2081 => x"b8",
          2082 => x"df",
          2083 => x"0b",
          2084 => x"33",
          2085 => x"06",
          2086 => x"82",
          2087 => x"06",
          2088 => x"91",
          2089 => x"f4",
          2090 => x"c3",
          2091 => x"0b",
          2092 => x"d8",
          2093 => x"c4",
          2094 => x"52",
          2095 => x"c3",
          2096 => x"5a",
          2097 => x"b7",
          2098 => x"7c",
          2099 => x"85",
          2100 => x"78",
          2101 => x"fd",
          2102 => x"10",
          2103 => x"c4",
          2104 => x"08",
          2105 => x"83",
          2106 => x"7e",
          2107 => x"3f",
          2108 => x"52",
          2109 => x"51",
          2110 => x"3f",
          2111 => x"08",
          2112 => x"81",
          2113 => x"38",
          2114 => x"3d",
          2115 => x"fb",
          2116 => x"d5",
          2117 => x"db",
          2118 => x"81",
          2119 => x"fe",
          2120 => x"d5",
          2121 => x"55",
          2122 => x"54",
          2123 => x"d5",
          2124 => x"51",
          2125 => x"fd",
          2126 => x"8c",
          2127 => x"ff",
          2128 => x"3f",
          2129 => x"81",
          2130 => x"bf",
          2131 => x"ef",
          2132 => x"c5",
          2133 => x"39",
          2134 => x"51",
          2135 => x"80",
          2136 => x"83",
          2137 => x"de",
          2138 => x"fd",
          2139 => x"39",
          2140 => x"84",
          2141 => x"80",
          2142 => x"8a",
          2143 => x"e4",
          2144 => x"fa",
          2145 => x"52",
          2146 => x"51",
          2147 => x"68",
          2148 => x"84",
          2149 => x"80",
          2150 => x"38",
          2151 => x"08",
          2152 => x"8c",
          2153 => x"3f",
          2154 => x"b8",
          2155 => x"11",
          2156 => x"05",
          2157 => x"3f",
          2158 => x"08",
          2159 => x"ff",
          2160 => x"83",
          2161 => x"d0",
          2162 => x"59",
          2163 => x"3d",
          2164 => x"53",
          2165 => x"51",
          2166 => x"84",
          2167 => x"80",
          2168 => x"38",
          2169 => x"f0",
          2170 => x"80",
          2171 => x"92",
          2172 => x"e4",
          2173 => x"38",
          2174 => x"08",
          2175 => x"83",
          2176 => x"d0",
          2177 => x"d4",
          2178 => x"80",
          2179 => x"51",
          2180 => x"7e",
          2181 => x"59",
          2182 => x"f9",
          2183 => x"9f",
          2184 => x"38",
          2185 => x"70",
          2186 => x"39",
          2187 => x"f4",
          2188 => x"80",
          2189 => x"ca",
          2190 => x"e4",
          2191 => x"f8",
          2192 => x"3d",
          2193 => x"53",
          2194 => x"51",
          2195 => x"84",
          2196 => x"86",
          2197 => x"59",
          2198 => x"78",
          2199 => x"d4",
          2200 => x"3f",
          2201 => x"08",
          2202 => x"52",
          2203 => x"b3",
          2204 => x"7e",
          2205 => x"ae",
          2206 => x"38",
          2207 => x"87",
          2208 => x"82",
          2209 => x"59",
          2210 => x"3d",
          2211 => x"53",
          2212 => x"51",
          2213 => x"84",
          2214 => x"80",
          2215 => x"38",
          2216 => x"fc",
          2217 => x"80",
          2218 => x"da",
          2219 => x"e4",
          2220 => x"f8",
          2221 => x"3d",
          2222 => x"53",
          2223 => x"51",
          2224 => x"84",
          2225 => x"80",
          2226 => x"38",
          2227 => x"51",
          2228 => x"68",
          2229 => x"78",
          2230 => x"8d",
          2231 => x"33",
          2232 => x"5c",
          2233 => x"2e",
          2234 => x"55",
          2235 => x"33",
          2236 => x"83",
          2237 => x"ce",
          2238 => x"66",
          2239 => x"19",
          2240 => x"59",
          2241 => x"3d",
          2242 => x"53",
          2243 => x"51",
          2244 => x"84",
          2245 => x"80",
          2246 => x"38",
          2247 => x"fc",
          2248 => x"80",
          2249 => x"de",
          2250 => x"e4",
          2251 => x"f7",
          2252 => x"3d",
          2253 => x"53",
          2254 => x"51",
          2255 => x"84",
          2256 => x"80",
          2257 => x"38",
          2258 => x"51",
          2259 => x"68",
          2260 => x"27",
          2261 => x"65",
          2262 => x"81",
          2263 => x"7c",
          2264 => x"05",
          2265 => x"b8",
          2266 => x"11",
          2267 => x"05",
          2268 => x"3f",
          2269 => x"08",
          2270 => x"c3",
          2271 => x"fe",
          2272 => x"ff",
          2273 => x"e7",
          2274 => x"b8",
          2275 => x"38",
          2276 => x"54",
          2277 => x"98",
          2278 => x"3f",
          2279 => x"08",
          2280 => x"52",
          2281 => x"fb",
          2282 => x"7e",
          2283 => x"ae",
          2284 => x"38",
          2285 => x"84",
          2286 => x"81",
          2287 => x"39",
          2288 => x"80",
          2289 => x"79",
          2290 => x"05",
          2291 => x"fe",
          2292 => x"ff",
          2293 => x"e7",
          2294 => x"b8",
          2295 => x"2e",
          2296 => x"68",
          2297 => x"db",
          2298 => x"34",
          2299 => x"49",
          2300 => x"fc",
          2301 => x"80",
          2302 => x"8a",
          2303 => x"e4",
          2304 => x"38",
          2305 => x"b8",
          2306 => x"11",
          2307 => x"05",
          2308 => x"3f",
          2309 => x"08",
          2310 => x"a3",
          2311 => x"fe",
          2312 => x"ff",
          2313 => x"e6",
          2314 => x"b8",
          2315 => x"2e",
          2316 => x"b8",
          2317 => x"11",
          2318 => x"05",
          2319 => x"3f",
          2320 => x"08",
          2321 => x"b8",
          2322 => x"83",
          2323 => x"cb",
          2324 => x"67",
          2325 => x"7a",
          2326 => x"65",
          2327 => x"70",
          2328 => x"0c",
          2329 => x"f5",
          2330 => x"d9",
          2331 => x"cf",
          2332 => x"ff",
          2333 => x"87",
          2334 => x"b8",
          2335 => x"3d",
          2336 => x"52",
          2337 => x"3f",
          2338 => x"b8",
          2339 => x"78",
          2340 => x"3f",
          2341 => x"08",
          2342 => x"a3",
          2343 => x"e4",
          2344 => x"f6",
          2345 => x"39",
          2346 => x"84",
          2347 => x"80",
          2348 => x"d2",
          2349 => x"e4",
          2350 => x"83",
          2351 => x"5a",
          2352 => x"83",
          2353 => x"f1",
          2354 => x"b8",
          2355 => x"11",
          2356 => x"05",
          2357 => x"3f",
          2358 => x"08",
          2359 => x"f1",
          2360 => x"79",
          2361 => x"8a",
          2362 => x"a4",
          2363 => x"3d",
          2364 => x"53",
          2365 => x"51",
          2366 => x"84",
          2367 => x"80",
          2368 => x"80",
          2369 => x"7a",
          2370 => x"38",
          2371 => x"90",
          2372 => x"70",
          2373 => x"2a",
          2374 => x"5f",
          2375 => x"2e",
          2376 => x"a0",
          2377 => x"88",
          2378 => x"b4",
          2379 => x"3f",
          2380 => x"54",
          2381 => x"52",
          2382 => x"a8",
          2383 => x"c0",
          2384 => x"3f",
          2385 => x"64",
          2386 => x"59",
          2387 => x"45",
          2388 => x"f0",
          2389 => x"80",
          2390 => x"a6",
          2391 => x"e4",
          2392 => x"f2",
          2393 => x"64",
          2394 => x"64",
          2395 => x"b8",
          2396 => x"11",
          2397 => x"05",
          2398 => x"3f",
          2399 => x"08",
          2400 => x"bb",
          2401 => x"02",
          2402 => x"22",
          2403 => x"05",
          2404 => x"45",
          2405 => x"f0",
          2406 => x"80",
          2407 => x"e2",
          2408 => x"e4",
          2409 => x"f2",
          2410 => x"5e",
          2411 => x"05",
          2412 => x"82",
          2413 => x"7d",
          2414 => x"fe",
          2415 => x"ff",
          2416 => x"e1",
          2417 => x"b8",
          2418 => x"b9",
          2419 => x"39",
          2420 => x"fc",
          2421 => x"80",
          2422 => x"aa",
          2423 => x"e4",
          2424 => x"81",
          2425 => x"5c",
          2426 => x"05",
          2427 => x"68",
          2428 => x"fb",
          2429 => x"3d",
          2430 => x"53",
          2431 => x"51",
          2432 => x"84",
          2433 => x"80",
          2434 => x"38",
          2435 => x"0c",
          2436 => x"05",
          2437 => x"f7",
          2438 => x"83",
          2439 => x"06",
          2440 => x"7b",
          2441 => x"ac",
          2442 => x"83",
          2443 => x"7c",
          2444 => x"3f",
          2445 => x"7b",
          2446 => x"da",
          2447 => x"8c",
          2448 => x"d8",
          2449 => x"3f",
          2450 => x"b8",
          2451 => x"11",
          2452 => x"05",
          2453 => x"3f",
          2454 => x"08",
          2455 => x"38",
          2456 => x"80",
          2457 => x"79",
          2458 => x"5b",
          2459 => x"f7",
          2460 => x"f1",
          2461 => x"7b",
          2462 => x"cf",
          2463 => x"ac",
          2464 => x"ea",
          2465 => x"e9",
          2466 => x"80",
          2467 => x"83",
          2468 => x"49",
          2469 => x"83",
          2470 => x"d3",
          2471 => x"59",
          2472 => x"83",
          2473 => x"d3",
          2474 => x"59",
          2475 => x"83",
          2476 => x"59",
          2477 => x"a5",
          2478 => x"b0",
          2479 => x"8b",
          2480 => x"84",
          2481 => x"3f",
          2482 => x"83",
          2483 => x"59",
          2484 => x"9b",
          2485 => x"b4",
          2486 => x"92",
          2487 => x"eb",
          2488 => x"80",
          2489 => x"83",
          2490 => x"49",
          2491 => x"83",
          2492 => x"5e",
          2493 => x"9b",
          2494 => x"bc",
          2495 => x"ee",
          2496 => x"e6",
          2497 => x"80",
          2498 => x"83",
          2499 => x"49",
          2500 => x"83",
          2501 => x"5d",
          2502 => x"94",
          2503 => x"c4",
          2504 => x"ca",
          2505 => x"d0",
          2506 => x"05",
          2507 => x"39",
          2508 => x"08",
          2509 => x"fb",
          2510 => x"3d",
          2511 => x"84",
          2512 => x"87",
          2513 => x"70",
          2514 => x"87",
          2515 => x"74",
          2516 => x"3f",
          2517 => x"08",
          2518 => x"08",
          2519 => x"84",
          2520 => x"51",
          2521 => x"74",
          2522 => x"08",
          2523 => x"87",
          2524 => x"70",
          2525 => x"87",
          2526 => x"74",
          2527 => x"3f",
          2528 => x"08",
          2529 => x"08",
          2530 => x"84",
          2531 => x"51",
          2532 => x"74",
          2533 => x"08",
          2534 => x"8c",
          2535 => x"87",
          2536 => x"0c",
          2537 => x"0b",
          2538 => x"94",
          2539 => x"e1",
          2540 => x"e0",
          2541 => x"84",
          2542 => x"34",
          2543 => x"d4",
          2544 => x"3d",
          2545 => x"0c",
          2546 => x"84",
          2547 => x"56",
          2548 => x"89",
          2549 => x"87",
          2550 => x"51",
          2551 => x"83",
          2552 => x"83",
          2553 => x"c4",
          2554 => x"f1",
          2555 => x"52",
          2556 => x"3f",
          2557 => x"54",
          2558 => x"53",
          2559 => x"52",
          2560 => x"51",
          2561 => x"8d",
          2562 => x"82",
          2563 => x"fb",
          2564 => x"70",
          2565 => x"80",
          2566 => x"74",
          2567 => x"83",
          2568 => x"70",
          2569 => x"52",
          2570 => x"2e",
          2571 => x"91",
          2572 => x"70",
          2573 => x"ff",
          2574 => x"55",
          2575 => x"f1",
          2576 => x"ff",
          2577 => x"a2",
          2578 => x"38",
          2579 => x"81",
          2580 => x"38",
          2581 => x"70",
          2582 => x"53",
          2583 => x"a0",
          2584 => x"81",
          2585 => x"2e",
          2586 => x"80",
          2587 => x"81",
          2588 => x"39",
          2589 => x"ff",
          2590 => x"70",
          2591 => x"81",
          2592 => x"81",
          2593 => x"32",
          2594 => x"80",
          2595 => x"52",
          2596 => x"80",
          2597 => x"80",
          2598 => x"05",
          2599 => x"76",
          2600 => x"70",
          2601 => x"0c",
          2602 => x"04",
          2603 => x"c4",
          2604 => x"2e",
          2605 => x"81",
          2606 => x"72",
          2607 => x"ff",
          2608 => x"54",
          2609 => x"e4",
          2610 => x"e0",
          2611 => x"55",
          2612 => x"53",
          2613 => x"09",
          2614 => x"f8",
          2615 => x"fc",
          2616 => x"53",
          2617 => x"38",
          2618 => x"b8",
          2619 => x"3d",
          2620 => x"3d",
          2621 => x"72",
          2622 => x"3f",
          2623 => x"08",
          2624 => x"38",
          2625 => x"e4",
          2626 => x"0d",
          2627 => x"0d",
          2628 => x"33",
          2629 => x"53",
          2630 => x"8b",
          2631 => x"38",
          2632 => x"ff",
          2633 => x"52",
          2634 => x"81",
          2635 => x"13",
          2636 => x"52",
          2637 => x"80",
          2638 => x"13",
          2639 => x"52",
          2640 => x"80",
          2641 => x"13",
          2642 => x"52",
          2643 => x"80",
          2644 => x"13",
          2645 => x"52",
          2646 => x"26",
          2647 => x"8a",
          2648 => x"87",
          2649 => x"e7",
          2650 => x"38",
          2651 => x"c0",
          2652 => x"72",
          2653 => x"98",
          2654 => x"13",
          2655 => x"98",
          2656 => x"13",
          2657 => x"98",
          2658 => x"13",
          2659 => x"98",
          2660 => x"13",
          2661 => x"98",
          2662 => x"13",
          2663 => x"98",
          2664 => x"87",
          2665 => x"0c",
          2666 => x"98",
          2667 => x"0b",
          2668 => x"9c",
          2669 => x"71",
          2670 => x"0c",
          2671 => x"04",
          2672 => x"7f",
          2673 => x"98",
          2674 => x"7d",
          2675 => x"98",
          2676 => x"7d",
          2677 => x"c0",
          2678 => x"5c",
          2679 => x"34",
          2680 => x"b4",
          2681 => x"83",
          2682 => x"c0",
          2683 => x"5c",
          2684 => x"34",
          2685 => x"ac",
          2686 => x"85",
          2687 => x"c0",
          2688 => x"5c",
          2689 => x"34",
          2690 => x"a4",
          2691 => x"88",
          2692 => x"c0",
          2693 => x"5a",
          2694 => x"23",
          2695 => x"79",
          2696 => x"06",
          2697 => x"ff",
          2698 => x"86",
          2699 => x"85",
          2700 => x"84",
          2701 => x"83",
          2702 => x"82",
          2703 => x"7d",
          2704 => x"06",
          2705 => x"88",
          2706 => x"bc",
          2707 => x"0d",
          2708 => x"0d",
          2709 => x"33",
          2710 => x"2e",
          2711 => x"51",
          2712 => x"3f",
          2713 => x"08",
          2714 => x"98",
          2715 => x"71",
          2716 => x"81",
          2717 => x"72",
          2718 => x"38",
          2719 => x"e4",
          2720 => x"0d",
          2721 => x"80",
          2722 => x"84",
          2723 => x"98",
          2724 => x"2c",
          2725 => x"ff",
          2726 => x"06",
          2727 => x"51",
          2728 => x"3f",
          2729 => x"08",
          2730 => x"98",
          2731 => x"71",
          2732 => x"38",
          2733 => x"3d",
          2734 => x"54",
          2735 => x"2b",
          2736 => x"80",
          2737 => x"84",
          2738 => x"98",
          2739 => x"2c",
          2740 => x"ff",
          2741 => x"73",
          2742 => x"14",
          2743 => x"73",
          2744 => x"71",
          2745 => x"0c",
          2746 => x"04",
          2747 => x"02",
          2748 => x"83",
          2749 => x"70",
          2750 => x"53",
          2751 => x"80",
          2752 => x"38",
          2753 => x"94",
          2754 => x"2a",
          2755 => x"53",
          2756 => x"80",
          2757 => x"71",
          2758 => x"81",
          2759 => x"70",
          2760 => x"81",
          2761 => x"53",
          2762 => x"8a",
          2763 => x"2a",
          2764 => x"71",
          2765 => x"81",
          2766 => x"87",
          2767 => x"52",
          2768 => x"86",
          2769 => x"94",
          2770 => x"72",
          2771 => x"b8",
          2772 => x"3d",
          2773 => x"91",
          2774 => x"06",
          2775 => x"97",
          2776 => x"32",
          2777 => x"72",
          2778 => x"38",
          2779 => x"81",
          2780 => x"80",
          2781 => x"87",
          2782 => x"08",
          2783 => x"70",
          2784 => x"54",
          2785 => x"38",
          2786 => x"3d",
          2787 => x"05",
          2788 => x"70",
          2789 => x"52",
          2790 => x"f1",
          2791 => x"3d",
          2792 => x"3d",
          2793 => x"80",
          2794 => x"56",
          2795 => x"77",
          2796 => x"38",
          2797 => x"f1",
          2798 => x"81",
          2799 => x"57",
          2800 => x"2e",
          2801 => x"87",
          2802 => x"08",
          2803 => x"70",
          2804 => x"54",
          2805 => x"2e",
          2806 => x"91",
          2807 => x"06",
          2808 => x"e3",
          2809 => x"32",
          2810 => x"72",
          2811 => x"38",
          2812 => x"81",
          2813 => x"cf",
          2814 => x"ff",
          2815 => x"c0",
          2816 => x"70",
          2817 => x"38",
          2818 => x"90",
          2819 => x"0c",
          2820 => x"33",
          2821 => x"ff",
          2822 => x"84",
          2823 => x"88",
          2824 => x"71",
          2825 => x"81",
          2826 => x"70",
          2827 => x"81",
          2828 => x"53",
          2829 => x"c1",
          2830 => x"2a",
          2831 => x"71",
          2832 => x"b5",
          2833 => x"94",
          2834 => x"96",
          2835 => x"06",
          2836 => x"70",
          2837 => x"39",
          2838 => x"87",
          2839 => x"08",
          2840 => x"8a",
          2841 => x"70",
          2842 => x"ab",
          2843 => x"9e",
          2844 => x"f1",
          2845 => x"c0",
          2846 => x"83",
          2847 => x"87",
          2848 => x"08",
          2849 => x"0c",
          2850 => x"98",
          2851 => x"ac",
          2852 => x"9e",
          2853 => x"f1",
          2854 => x"c0",
          2855 => x"83",
          2856 => x"87",
          2857 => x"08",
          2858 => x"0c",
          2859 => x"b0",
          2860 => x"bc",
          2861 => x"9e",
          2862 => x"f1",
          2863 => x"c0",
          2864 => x"83",
          2865 => x"87",
          2866 => x"08",
          2867 => x"0c",
          2868 => x"c0",
          2869 => x"cc",
          2870 => x"9e",
          2871 => x"f1",
          2872 => x"c0",
          2873 => x"52",
          2874 => x"d4",
          2875 => x"9e",
          2876 => x"f1",
          2877 => x"c0",
          2878 => x"83",
          2879 => x"87",
          2880 => x"08",
          2881 => x"0c",
          2882 => x"f1",
          2883 => x"0b",
          2884 => x"90",
          2885 => x"80",
          2886 => x"52",
          2887 => x"fb",
          2888 => x"f1",
          2889 => x"0b",
          2890 => x"90",
          2891 => x"80",
          2892 => x"52",
          2893 => x"2e",
          2894 => x"52",
          2895 => x"e6",
          2896 => x"87",
          2897 => x"08",
          2898 => x"0a",
          2899 => x"52",
          2900 => x"83",
          2901 => x"71",
          2902 => x"34",
          2903 => x"c0",
          2904 => x"70",
          2905 => x"06",
          2906 => x"70",
          2907 => x"38",
          2908 => x"83",
          2909 => x"80",
          2910 => x"9e",
          2911 => x"a0",
          2912 => x"51",
          2913 => x"80",
          2914 => x"81",
          2915 => x"f1",
          2916 => x"0b",
          2917 => x"90",
          2918 => x"80",
          2919 => x"52",
          2920 => x"2e",
          2921 => x"52",
          2922 => x"ea",
          2923 => x"87",
          2924 => x"08",
          2925 => x"80",
          2926 => x"52",
          2927 => x"83",
          2928 => x"71",
          2929 => x"34",
          2930 => x"c0",
          2931 => x"70",
          2932 => x"06",
          2933 => x"70",
          2934 => x"38",
          2935 => x"83",
          2936 => x"80",
          2937 => x"9e",
          2938 => x"81",
          2939 => x"51",
          2940 => x"80",
          2941 => x"81",
          2942 => x"f1",
          2943 => x"0b",
          2944 => x"90",
          2945 => x"c0",
          2946 => x"52",
          2947 => x"2e",
          2948 => x"52",
          2949 => x"ee",
          2950 => x"87",
          2951 => x"08",
          2952 => x"06",
          2953 => x"70",
          2954 => x"38",
          2955 => x"83",
          2956 => x"87",
          2957 => x"08",
          2958 => x"70",
          2959 => x"51",
          2960 => x"f0",
          2961 => x"87",
          2962 => x"08",
          2963 => x"06",
          2964 => x"70",
          2965 => x"38",
          2966 => x"83",
          2967 => x"87",
          2968 => x"08",
          2969 => x"70",
          2970 => x"51",
          2971 => x"f2",
          2972 => x"87",
          2973 => x"08",
          2974 => x"51",
          2975 => x"80",
          2976 => x"81",
          2977 => x"f1",
          2978 => x"c0",
          2979 => x"87",
          2980 => x"83",
          2981 => x"83",
          2982 => x"81",
          2983 => x"39",
          2984 => x"83",
          2985 => x"ff",
          2986 => x"83",
          2987 => x"54",
          2988 => x"38",
          2989 => x"51",
          2990 => x"83",
          2991 => x"55",
          2992 => x"38",
          2993 => x"33",
          2994 => x"d1",
          2995 => x"e8",
          2996 => x"85",
          2997 => x"f1",
          2998 => x"74",
          2999 => x"83",
          3000 => x"54",
          3001 => x"38",
          3002 => x"33",
          3003 => x"b3",
          3004 => x"f3",
          3005 => x"84",
          3006 => x"f1",
          3007 => x"74",
          3008 => x"83",
          3009 => x"56",
          3010 => x"38",
          3011 => x"33",
          3012 => x"b1",
          3013 => x"ec",
          3014 => x"83",
          3015 => x"f1",
          3016 => x"75",
          3017 => x"83",
          3018 => x"54",
          3019 => x"38",
          3020 => x"51",
          3021 => x"83",
          3022 => x"52",
          3023 => x"51",
          3024 => x"3f",
          3025 => x"08",
          3026 => x"80",
          3027 => x"b8",
          3028 => x"d0",
          3029 => x"d9",
          3030 => x"b5",
          3031 => x"d9",
          3032 => x"8f",
          3033 => x"d4",
          3034 => x"d9",
          3035 => x"b5",
          3036 => x"f1",
          3037 => x"bd",
          3038 => x"75",
          3039 => x"3f",
          3040 => x"08",
          3041 => x"29",
          3042 => x"54",
          3043 => x"e4",
          3044 => x"da",
          3045 => x"b4",
          3046 => x"f1",
          3047 => x"74",
          3048 => x"83",
          3049 => x"55",
          3050 => x"8a",
          3051 => x"3f",
          3052 => x"04",
          3053 => x"08",
          3054 => x"c0",
          3055 => x"c9",
          3056 => x"b8",
          3057 => x"84",
          3058 => x"71",
          3059 => x"84",
          3060 => x"52",
          3061 => x"51",
          3062 => x"3f",
          3063 => x"fe",
          3064 => x"0d",
          3065 => x"dc",
          3066 => x"84",
          3067 => x"51",
          3068 => x"84",
          3069 => x"bd",
          3070 => x"76",
          3071 => x"54",
          3072 => x"08",
          3073 => x"d8",
          3074 => x"fc",
          3075 => x"e6",
          3076 => x"80",
          3077 => x"38",
          3078 => x"83",
          3079 => x"c0",
          3080 => x"d8",
          3081 => x"cb",
          3082 => x"c8",
          3083 => x"d8",
          3084 => x"b3",
          3085 => x"f1",
          3086 => x"83",
          3087 => x"ff",
          3088 => x"83",
          3089 => x"52",
          3090 => x"51",
          3091 => x"3f",
          3092 => x"51",
          3093 => x"83",
          3094 => x"52",
          3095 => x"51",
          3096 => x"3f",
          3097 => x"08",
          3098 => x"c0",
          3099 => x"c8",
          3100 => x"b8",
          3101 => x"84",
          3102 => x"71",
          3103 => x"84",
          3104 => x"52",
          3105 => x"51",
          3106 => x"3f",
          3107 => x"33",
          3108 => x"2e",
          3109 => x"fe",
          3110 => x"db",
          3111 => x"bf",
          3112 => x"f1",
          3113 => x"73",
          3114 => x"84",
          3115 => x"39",
          3116 => x"51",
          3117 => x"3f",
          3118 => x"33",
          3119 => x"2e",
          3120 => x"d6",
          3121 => x"a0",
          3122 => x"a7",
          3123 => x"ec",
          3124 => x"80",
          3125 => x"38",
          3126 => x"db",
          3127 => x"bf",
          3128 => x"f1",
          3129 => x"73",
          3130 => x"a9",
          3131 => x"83",
          3132 => x"52",
          3133 => x"51",
          3134 => x"3f",
          3135 => x"33",
          3136 => x"2e",
          3137 => x"d2",
          3138 => x"f4",
          3139 => x"db",
          3140 => x"b1",
          3141 => x"f1",
          3142 => x"74",
          3143 => x"e3",
          3144 => x"83",
          3145 => x"52",
          3146 => x"51",
          3147 => x"3f",
          3148 => x"33",
          3149 => x"2e",
          3150 => x"cd",
          3151 => x"b0",
          3152 => x"b4",
          3153 => x"52",
          3154 => x"51",
          3155 => x"3f",
          3156 => x"33",
          3157 => x"2e",
          3158 => x"c7",
          3159 => x"a8",
          3160 => x"ac",
          3161 => x"52",
          3162 => x"51",
          3163 => x"3f",
          3164 => x"33",
          3165 => x"2e",
          3166 => x"c1",
          3167 => x"a0",
          3168 => x"a4",
          3169 => x"52",
          3170 => x"51",
          3171 => x"3f",
          3172 => x"33",
          3173 => x"2e",
          3174 => x"c1",
          3175 => x"b8",
          3176 => x"bc",
          3177 => x"52",
          3178 => x"51",
          3179 => x"3f",
          3180 => x"33",
          3181 => x"2e",
          3182 => x"c1",
          3183 => x"c0",
          3184 => x"c4",
          3185 => x"52",
          3186 => x"51",
          3187 => x"3f",
          3188 => x"33",
          3189 => x"2e",
          3190 => x"c1",
          3191 => x"ac",
          3192 => x"a4",
          3193 => x"b4",
          3194 => x"87",
          3195 => x"e6",
          3196 => x"80",
          3197 => x"38",
          3198 => x"3d",
          3199 => x"05",
          3200 => x"85",
          3201 => x"71",
          3202 => x"c2",
          3203 => x"71",
          3204 => x"dd",
          3205 => x"af",
          3206 => x"3d",
          3207 => x"dd",
          3208 => x"af",
          3209 => x"3d",
          3210 => x"dd",
          3211 => x"af",
          3212 => x"3d",
          3213 => x"dd",
          3214 => x"af",
          3215 => x"3d",
          3216 => x"dd",
          3217 => x"af",
          3218 => x"3d",
          3219 => x"dd",
          3220 => x"af",
          3221 => x"3d",
          3222 => x"88",
          3223 => x"80",
          3224 => x"96",
          3225 => x"83",
          3226 => x"87",
          3227 => x"0c",
          3228 => x"0d",
          3229 => x"ad",
          3230 => x"5a",
          3231 => x"58",
          3232 => x"f2",
          3233 => x"82",
          3234 => x"84",
          3235 => x"80",
          3236 => x"3d",
          3237 => x"83",
          3238 => x"54",
          3239 => x"52",
          3240 => x"d2",
          3241 => x"b8",
          3242 => x"2e",
          3243 => x"51",
          3244 => x"84",
          3245 => x"81",
          3246 => x"80",
          3247 => x"e4",
          3248 => x"38",
          3249 => x"08",
          3250 => x"18",
          3251 => x"74",
          3252 => x"70",
          3253 => x"07",
          3254 => x"55",
          3255 => x"2e",
          3256 => x"ff",
          3257 => x"f2",
          3258 => x"11",
          3259 => x"82",
          3260 => x"84",
          3261 => x"8f",
          3262 => x"2e",
          3263 => x"84",
          3264 => x"a9",
          3265 => x"83",
          3266 => x"ff",
          3267 => x"78",
          3268 => x"81",
          3269 => x"76",
          3270 => x"c0",
          3271 => x"51",
          3272 => x"ab",
          3273 => x"84",
          3274 => x"76",
          3275 => x"83",
          3276 => x"ff",
          3277 => x"80",
          3278 => x"e4",
          3279 => x"0d",
          3280 => x"0d",
          3281 => x"ad",
          3282 => x"72",
          3283 => x"57",
          3284 => x"73",
          3285 => x"91",
          3286 => x"8d",
          3287 => x"75",
          3288 => x"83",
          3289 => x"70",
          3290 => x"ff",
          3291 => x"84",
          3292 => x"53",
          3293 => x"08",
          3294 => x"3f",
          3295 => x"08",
          3296 => x"14",
          3297 => x"81",
          3298 => x"38",
          3299 => x"99",
          3300 => x"70",
          3301 => x"57",
          3302 => x"27",
          3303 => x"54",
          3304 => x"e4",
          3305 => x"0d",
          3306 => x"5a",
          3307 => x"84",
          3308 => x"80",
          3309 => x"ce",
          3310 => x"e4",
          3311 => x"d1",
          3312 => x"53",
          3313 => x"51",
          3314 => x"84",
          3315 => x"81",
          3316 => x"73",
          3317 => x"38",
          3318 => x"81",
          3319 => x"54",
          3320 => x"fe",
          3321 => x"b6",
          3322 => x"77",
          3323 => x"76",
          3324 => x"38",
          3325 => x"5b",
          3326 => x"55",
          3327 => x"09",
          3328 => x"d5",
          3329 => x"26",
          3330 => x"0b",
          3331 => x"56",
          3332 => x"73",
          3333 => x"08",
          3334 => x"d0",
          3335 => x"82",
          3336 => x"84",
          3337 => x"80",
          3338 => x"f2",
          3339 => x"80",
          3340 => x"51",
          3341 => x"3f",
          3342 => x"08",
          3343 => x"38",
          3344 => x"bd",
          3345 => x"b8",
          3346 => x"80",
          3347 => x"e4",
          3348 => x"38",
          3349 => x"08",
          3350 => x"19",
          3351 => x"77",
          3352 => x"75",
          3353 => x"83",
          3354 => x"56",
          3355 => x"3f",
          3356 => x"09",
          3357 => x"b2",
          3358 => x"84",
          3359 => x"aa",
          3360 => x"ce",
          3361 => x"3d",
          3362 => x"08",
          3363 => x"5a",
          3364 => x"0b",
          3365 => x"83",
          3366 => x"83",
          3367 => x"56",
          3368 => x"38",
          3369 => x"cc",
          3370 => x"74",
          3371 => x"cb",
          3372 => x"2e",
          3373 => x"81",
          3374 => x"5a",
          3375 => x"a0",
          3376 => x"2e",
          3377 => x"93",
          3378 => x"5f",
          3379 => x"eb",
          3380 => x"b8",
          3381 => x"2b",
          3382 => x"5b",
          3383 => x"2e",
          3384 => x"81",
          3385 => x"d0",
          3386 => x"98",
          3387 => x"2c",
          3388 => x"33",
          3389 => x"70",
          3390 => x"98",
          3391 => x"10",
          3392 => x"ec",
          3393 => x"15",
          3394 => x"53",
          3395 => x"52",
          3396 => x"59",
          3397 => x"79",
          3398 => x"38",
          3399 => x"81",
          3400 => x"81",
          3401 => x"81",
          3402 => x"70",
          3403 => x"55",
          3404 => x"81",
          3405 => x"10",
          3406 => x"2b",
          3407 => x"0b",
          3408 => x"16",
          3409 => x"77",
          3410 => x"38",
          3411 => x"15",
          3412 => x"33",
          3413 => x"75",
          3414 => x"38",
          3415 => x"c2",
          3416 => x"d0",
          3417 => x"57",
          3418 => x"81",
          3419 => x"1b",
          3420 => x"70",
          3421 => x"d0",
          3422 => x"98",
          3423 => x"2c",
          3424 => x"05",
          3425 => x"83",
          3426 => x"33",
          3427 => x"5d",
          3428 => x"57",
          3429 => x"81",
          3430 => x"84",
          3431 => x"fe",
          3432 => x"57",
          3433 => x"38",
          3434 => x"0a",
          3435 => x"0a",
          3436 => x"2c",
          3437 => x"06",
          3438 => x"76",
          3439 => x"c0",
          3440 => x"16",
          3441 => x"51",
          3442 => x"83",
          3443 => x"33",
          3444 => x"61",
          3445 => x"83",
          3446 => x"08",
          3447 => x"42",
          3448 => x"2e",
          3449 => x"76",
          3450 => x"bc",
          3451 => x"39",
          3452 => x"80",
          3453 => x"38",
          3454 => x"81",
          3455 => x"39",
          3456 => x"fe",
          3457 => x"84",
          3458 => x"76",
          3459 => x"34",
          3460 => x"76",
          3461 => x"55",
          3462 => x"fd",
          3463 => x"10",
          3464 => x"84",
          3465 => x"08",
          3466 => x"f4",
          3467 => x"0c",
          3468 => x"d0",
          3469 => x"0b",
          3470 => x"34",
          3471 => x"d0",
          3472 => x"75",
          3473 => x"85",
          3474 => x"c8",
          3475 => x"51",
          3476 => x"3f",
          3477 => x"33",
          3478 => x"76",
          3479 => x"34",
          3480 => x"84",
          3481 => x"70",
          3482 => x"84",
          3483 => x"5b",
          3484 => x"79",
          3485 => x"38",
          3486 => x"08",
          3487 => x"58",
          3488 => x"a8",
          3489 => x"70",
          3490 => x"ff",
          3491 => x"fc",
          3492 => x"93",
          3493 => x"38",
          3494 => x"83",
          3495 => x"70",
          3496 => x"75",
          3497 => x"75",
          3498 => x"34",
          3499 => x"84",
          3500 => x"84",
          3501 => x"56",
          3502 => x"2e",
          3503 => x"d4",
          3504 => x"88",
          3505 => x"a6",
          3506 => x"c8",
          3507 => x"51",
          3508 => x"3f",
          3509 => x"08",
          3510 => x"ff",
          3511 => x"84",
          3512 => x"ff",
          3513 => x"84",
          3514 => x"7a",
          3515 => x"55",
          3516 => x"7b",
          3517 => x"90",
          3518 => x"d0",
          3519 => x"cd",
          3520 => x"38",
          3521 => x"08",
          3522 => x"9e",
          3523 => x"10",
          3524 => x"05",
          3525 => x"57",
          3526 => x"f9",
          3527 => x"56",
          3528 => x"fb",
          3529 => x"51",
          3530 => x"3f",
          3531 => x"08",
          3532 => x"34",
          3533 => x"08",
          3534 => x"81",
          3535 => x"52",
          3536 => x"b8",
          3537 => x"d0",
          3538 => x"d0",
          3539 => x"56",
          3540 => x"ff",
          3541 => x"d4",
          3542 => x"88",
          3543 => x"8e",
          3544 => x"c8",
          3545 => x"51",
          3546 => x"3f",
          3547 => x"08",
          3548 => x"ff",
          3549 => x"84",
          3550 => x"ff",
          3551 => x"84",
          3552 => x"74",
          3553 => x"55",
          3554 => x"d0",
          3555 => x"81",
          3556 => x"d0",
          3557 => x"57",
          3558 => x"27",
          3559 => x"84",
          3560 => x"52",
          3561 => x"76",
          3562 => x"34",
          3563 => x"33",
          3564 => x"b3",
          3565 => x"d0",
          3566 => x"81",
          3567 => x"d0",
          3568 => x"57",
          3569 => x"27",
          3570 => x"84",
          3571 => x"52",
          3572 => x"76",
          3573 => x"34",
          3574 => x"33",
          3575 => x"b3",
          3576 => x"d0",
          3577 => x"81",
          3578 => x"d0",
          3579 => x"57",
          3580 => x"26",
          3581 => x"f9",
          3582 => x"d0",
          3583 => x"d0",
          3584 => x"56",
          3585 => x"f9",
          3586 => x"15",
          3587 => x"d0",
          3588 => x"98",
          3589 => x"2c",
          3590 => x"06",
          3591 => x"60",
          3592 => x"ef",
          3593 => x"c8",
          3594 => x"51",
          3595 => x"3f",
          3596 => x"33",
          3597 => x"70",
          3598 => x"d0",
          3599 => x"57",
          3600 => x"77",
          3601 => x"38",
          3602 => x"08",
          3603 => x"ff",
          3604 => x"74",
          3605 => x"29",
          3606 => x"05",
          3607 => x"84",
          3608 => x"5d",
          3609 => x"7b",
          3610 => x"38",
          3611 => x"08",
          3612 => x"ff",
          3613 => x"74",
          3614 => x"29",
          3615 => x"05",
          3616 => x"84",
          3617 => x"5d",
          3618 => x"75",
          3619 => x"38",
          3620 => x"7b",
          3621 => x"18",
          3622 => x"84",
          3623 => x"52",
          3624 => x"ff",
          3625 => x"75",
          3626 => x"29",
          3627 => x"05",
          3628 => x"84",
          3629 => x"5b",
          3630 => x"79",
          3631 => x"38",
          3632 => x"81",
          3633 => x"34",
          3634 => x"08",
          3635 => x"51",
          3636 => x"3f",
          3637 => x"0a",
          3638 => x"0a",
          3639 => x"2c",
          3640 => x"33",
          3641 => x"78",
          3642 => x"a7",
          3643 => x"39",
          3644 => x"33",
          3645 => x"2e",
          3646 => x"84",
          3647 => x"52",
          3648 => x"b0",
          3649 => x"d0",
          3650 => x"05",
          3651 => x"d0",
          3652 => x"81",
          3653 => x"dd",
          3654 => x"a4",
          3655 => x"5f",
          3656 => x"84",
          3657 => x"52",
          3658 => x"b0",
          3659 => x"d0",
          3660 => x"51",
          3661 => x"84",
          3662 => x"81",
          3663 => x"77",
          3664 => x"84",
          3665 => x"57",
          3666 => x"80",
          3667 => x"f2",
          3668 => x"10",
          3669 => x"fc",
          3670 => x"57",
          3671 => x"8b",
          3672 => x"82",
          3673 => x"06",
          3674 => x"05",
          3675 => x"53",
          3676 => x"e7",
          3677 => x"b8",
          3678 => x"0c",
          3679 => x"33",
          3680 => x"83",
          3681 => x"70",
          3682 => x"41",
          3683 => x"38",
          3684 => x"08",
          3685 => x"2e",
          3686 => x"f2",
          3687 => x"77",
          3688 => x"bc",
          3689 => x"84",
          3690 => x"80",
          3691 => x"a4",
          3692 => x"b8",
          3693 => x"3d",
          3694 => x"d0",
          3695 => x"74",
          3696 => x"38",
          3697 => x"08",
          3698 => x"ff",
          3699 => x"84",
          3700 => x"52",
          3701 => x"af",
          3702 => x"d4",
          3703 => x"88",
          3704 => x"8a",
          3705 => x"a8",
          3706 => x"56",
          3707 => x"a8",
          3708 => x"ff",
          3709 => x"cc",
          3710 => x"e0",
          3711 => x"88",
          3712 => x"84",
          3713 => x"80",
          3714 => x"a4",
          3715 => x"39",
          3716 => x"80",
          3717 => x"34",
          3718 => x"33",
          3719 => x"2e",
          3720 => x"d4",
          3721 => x"88",
          3722 => x"c2",
          3723 => x"c8",
          3724 => x"51",
          3725 => x"3f",
          3726 => x"08",
          3727 => x"ff",
          3728 => x"84",
          3729 => x"ff",
          3730 => x"84",
          3731 => x"7c",
          3732 => x"55",
          3733 => x"83",
          3734 => x"ff",
          3735 => x"80",
          3736 => x"a8",
          3737 => x"84",
          3738 => x"7b",
          3739 => x"0c",
          3740 => x"04",
          3741 => x"33",
          3742 => x"06",
          3743 => x"80",
          3744 => x"38",
          3745 => x"33",
          3746 => x"78",
          3747 => x"34",
          3748 => x"77",
          3749 => x"34",
          3750 => x"08",
          3751 => x"ff",
          3752 => x"84",
          3753 => x"70",
          3754 => x"98",
          3755 => x"a4",
          3756 => x"5b",
          3757 => x"24",
          3758 => x"84",
          3759 => x"52",
          3760 => x"ad",
          3761 => x"d0",
          3762 => x"98",
          3763 => x"2c",
          3764 => x"33",
          3765 => x"56",
          3766 => x"f3",
          3767 => x"d4",
          3768 => x"88",
          3769 => x"86",
          3770 => x"80",
          3771 => x"80",
          3772 => x"98",
          3773 => x"a4",
          3774 => x"55",
          3775 => x"f3",
          3776 => x"d4",
          3777 => x"88",
          3778 => x"e2",
          3779 => x"80",
          3780 => x"80",
          3781 => x"98",
          3782 => x"a4",
          3783 => x"55",
          3784 => x"ff",
          3785 => x"a5",
          3786 => x"57",
          3787 => x"77",
          3788 => x"c8",
          3789 => x"33",
          3790 => x"b2",
          3791 => x"80",
          3792 => x"80",
          3793 => x"98",
          3794 => x"a4",
          3795 => x"5b",
          3796 => x"fe",
          3797 => x"16",
          3798 => x"33",
          3799 => x"d4",
          3800 => x"76",
          3801 => x"ac",
          3802 => x"81",
          3803 => x"81",
          3804 => x"70",
          3805 => x"d0",
          3806 => x"57",
          3807 => x"24",
          3808 => x"fe",
          3809 => x"d0",
          3810 => x"81",
          3811 => x"58",
          3812 => x"f2",
          3813 => x"d0",
          3814 => x"76",
          3815 => x"38",
          3816 => x"70",
          3817 => x"41",
          3818 => x"a1",
          3819 => x"5b",
          3820 => x"1c",
          3821 => x"80",
          3822 => x"ff",
          3823 => x"98",
          3824 => x"a8",
          3825 => x"58",
          3826 => x"e1",
          3827 => x"55",
          3828 => x"a8",
          3829 => x"ff",
          3830 => x"5a",
          3831 => x"7a",
          3832 => x"a4",
          3833 => x"60",
          3834 => x"81",
          3835 => x"84",
          3836 => x"75",
          3837 => x"a8",
          3838 => x"80",
          3839 => x"ff",
          3840 => x"98",
          3841 => x"ff",
          3842 => x"5c",
          3843 => x"24",
          3844 => x"77",
          3845 => x"98",
          3846 => x"ff",
          3847 => x"59",
          3848 => x"f1",
          3849 => x"d4",
          3850 => x"88",
          3851 => x"be",
          3852 => x"80",
          3853 => x"80",
          3854 => x"98",
          3855 => x"a4",
          3856 => x"41",
          3857 => x"f1",
          3858 => x"d4",
          3859 => x"88",
          3860 => x"9a",
          3861 => x"80",
          3862 => x"80",
          3863 => x"98",
          3864 => x"a4",
          3865 => x"41",
          3866 => x"ff",
          3867 => x"dd",
          3868 => x"fc",
          3869 => x"80",
          3870 => x"38",
          3871 => x"ad",
          3872 => x"b8",
          3873 => x"d0",
          3874 => x"b8",
          3875 => x"ff",
          3876 => x"53",
          3877 => x"51",
          3878 => x"3f",
          3879 => x"33",
          3880 => x"33",
          3881 => x"80",
          3882 => x"38",
          3883 => x"08",
          3884 => x"ff",
          3885 => x"84",
          3886 => x"52",
          3887 => x"a9",
          3888 => x"d4",
          3889 => x"88",
          3890 => x"a2",
          3891 => x"a8",
          3892 => x"5b",
          3893 => x"a8",
          3894 => x"ff",
          3895 => x"39",
          3896 => x"e1",
          3897 => x"b8",
          3898 => x"f2",
          3899 => x"b8",
          3900 => x"a5",
          3901 => x"f2",
          3902 => x"ef",
          3903 => x"c3",
          3904 => x"c8",
          3905 => x"16",
          3906 => x"58",
          3907 => x"3f",
          3908 => x"0a",
          3909 => x"0a",
          3910 => x"2c",
          3911 => x"33",
          3912 => x"76",
          3913 => x"38",
          3914 => x"33",
          3915 => x"70",
          3916 => x"81",
          3917 => x"58",
          3918 => x"7a",
          3919 => x"38",
          3920 => x"83",
          3921 => x"80",
          3922 => x"38",
          3923 => x"57",
          3924 => x"08",
          3925 => x"38",
          3926 => x"18",
          3927 => x"80",
          3928 => x"80",
          3929 => x"d4",
          3930 => x"d0",
          3931 => x"80",
          3932 => x"38",
          3933 => x"e7",
          3934 => x"f2",
          3935 => x"80",
          3936 => x"80",
          3937 => x"d0",
          3938 => x"b4",
          3939 => x"ee",
          3940 => x"51",
          3941 => x"3f",
          3942 => x"ff",
          3943 => x"58",
          3944 => x"25",
          3945 => x"ff",
          3946 => x"51",
          3947 => x"3f",
          3948 => x"08",
          3949 => x"34",
          3950 => x"08",
          3951 => x"81",
          3952 => x"52",
          3953 => x"ab",
          3954 => x"0b",
          3955 => x"33",
          3956 => x"33",
          3957 => x"74",
          3958 => x"97",
          3959 => x"c8",
          3960 => x"51",
          3961 => x"3f",
          3962 => x"08",
          3963 => x"ff",
          3964 => x"84",
          3965 => x"52",
          3966 => x"a6",
          3967 => x"d0",
          3968 => x"05",
          3969 => x"d0",
          3970 => x"81",
          3971 => x"c7",
          3972 => x"34",
          3973 => x"d0",
          3974 => x"0b",
          3975 => x"34",
          3976 => x"e4",
          3977 => x"0d",
          3978 => x"ff",
          3979 => x"84",
          3980 => x"84",
          3981 => x"84",
          3982 => x"81",
          3983 => x"05",
          3984 => x"7b",
          3985 => x"a2",
          3986 => x"70",
          3987 => x"84",
          3988 => x"84",
          3989 => x"58",
          3990 => x"74",
          3991 => x"93",
          3992 => x"c8",
          3993 => x"51",
          3994 => x"3f",
          3995 => x"08",
          3996 => x"ff",
          3997 => x"84",
          3998 => x"52",
          3999 => x"a5",
          4000 => x"d0",
          4001 => x"05",
          4002 => x"d0",
          4003 => x"81",
          4004 => x"c7",
          4005 => x"ff",
          4006 => x"84",
          4007 => x"84",
          4008 => x"84",
          4009 => x"81",
          4010 => x"05",
          4011 => x"7b",
          4012 => x"b6",
          4013 => x"70",
          4014 => x"84",
          4015 => x"84",
          4016 => x"58",
          4017 => x"74",
          4018 => x"a7",
          4019 => x"c8",
          4020 => x"51",
          4021 => x"3f",
          4022 => x"08",
          4023 => x"ff",
          4024 => x"84",
          4025 => x"52",
          4026 => x"a5",
          4027 => x"d0",
          4028 => x"05",
          4029 => x"d0",
          4030 => x"81",
          4031 => x"c7",
          4032 => x"80",
          4033 => x"83",
          4034 => x"70",
          4035 => x"fc",
          4036 => x"fc",
          4037 => x"70",
          4038 => x"56",
          4039 => x"3f",
          4040 => x"08",
          4041 => x"f2",
          4042 => x"10",
          4043 => x"fc",
          4044 => x"57",
          4045 => x"80",
          4046 => x"38",
          4047 => x"52",
          4048 => x"a8",
          4049 => x"f2",
          4050 => x"05",
          4051 => x"06",
          4052 => x"79",
          4053 => x"38",
          4054 => x"d4",
          4055 => x"39",
          4056 => x"f8",
          4057 => x"53",
          4058 => x"51",
          4059 => x"3f",
          4060 => x"08",
          4061 => x"82",
          4062 => x"83",
          4063 => x"51",
          4064 => x"3f",
          4065 => x"d0",
          4066 => x"0b",
          4067 => x"34",
          4068 => x"e4",
          4069 => x"0d",
          4070 => x"77",
          4071 => x"e4",
          4072 => x"c9",
          4073 => x"b8",
          4074 => x"a5",
          4075 => x"e4",
          4076 => x"5c",
          4077 => x"d0",
          4078 => x"f8",
          4079 => x"82",
          4080 => x"84",
          4081 => x"5a",
          4082 => x"08",
          4083 => x"81",
          4084 => x"38",
          4085 => x"08",
          4086 => x"cc",
          4087 => x"e4",
          4088 => x"0b",
          4089 => x"08",
          4090 => x"38",
          4091 => x"08",
          4092 => x"1b",
          4093 => x"77",
          4094 => x"ff",
          4095 => x"d4",
          4096 => x"10",
          4097 => x"05",
          4098 => x"40",
          4099 => x"80",
          4100 => x"82",
          4101 => x"06",
          4102 => x"05",
          4103 => x"53",
          4104 => x"da",
          4105 => x"b8",
          4106 => x"0c",
          4107 => x"33",
          4108 => x"83",
          4109 => x"70",
          4110 => x"41",
          4111 => x"81",
          4112 => x"ff",
          4113 => x"93",
          4114 => x"38",
          4115 => x"ff",
          4116 => x"06",
          4117 => x"77",
          4118 => x"f9",
          4119 => x"53",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"33",
          4123 => x"81",
          4124 => x"57",
          4125 => x"80",
          4126 => x"0b",
          4127 => x"34",
          4128 => x"74",
          4129 => x"f8",
          4130 => x"d4",
          4131 => x"2b",
          4132 => x"83",
          4133 => x"81",
          4134 => x"52",
          4135 => x"d9",
          4136 => x"b8",
          4137 => x"0c",
          4138 => x"33",
          4139 => x"83",
          4140 => x"70",
          4141 => x"41",
          4142 => x"ff",
          4143 => x"9e",
          4144 => x"f2",
          4145 => x"f7",
          4146 => x"f2",
          4147 => x"c0",
          4148 => x"cc",
          4149 => x"9b",
          4150 => x"eb",
          4151 => x"39",
          4152 => x"02",
          4153 => x"33",
          4154 => x"80",
          4155 => x"5b",
          4156 => x"26",
          4157 => x"72",
          4158 => x"8b",
          4159 => x"25",
          4160 => x"72",
          4161 => x"a8",
          4162 => x"a0",
          4163 => x"a7",
          4164 => x"5e",
          4165 => x"9f",
          4166 => x"76",
          4167 => x"75",
          4168 => x"34",
          4169 => x"95",
          4170 => x"f8",
          4171 => x"f8",
          4172 => x"98",
          4173 => x"2b",
          4174 => x"2b",
          4175 => x"7a",
          4176 => x"56",
          4177 => x"27",
          4178 => x"74",
          4179 => x"56",
          4180 => x"70",
          4181 => x"0c",
          4182 => x"ee",
          4183 => x"27",
          4184 => x"f8",
          4185 => x"97",
          4186 => x"78",
          4187 => x"55",
          4188 => x"e0",
          4189 => x"74",
          4190 => x"56",
          4191 => x"53",
          4192 => x"90",
          4193 => x"86",
          4194 => x"0b",
          4195 => x"33",
          4196 => x"11",
          4197 => x"33",
          4198 => x"11",
          4199 => x"41",
          4200 => x"86",
          4201 => x"0b",
          4202 => x"33",
          4203 => x"06",
          4204 => x"33",
          4205 => x"06",
          4206 => x"22",
          4207 => x"ff",
          4208 => x"29",
          4209 => x"58",
          4210 => x"5d",
          4211 => x"87",
          4212 => x"31",
          4213 => x"79",
          4214 => x"7e",
          4215 => x"7c",
          4216 => x"7a",
          4217 => x"06",
          4218 => x"06",
          4219 => x"14",
          4220 => x"57",
          4221 => x"74",
          4222 => x"83",
          4223 => x"74",
          4224 => x"70",
          4225 => x"59",
          4226 => x"06",
          4227 => x"2e",
          4228 => x"78",
          4229 => x"72",
          4230 => x"c1",
          4231 => x"70",
          4232 => x"34",
          4233 => x"33",
          4234 => x"05",
          4235 => x"39",
          4236 => x"80",
          4237 => x"b0",
          4238 => x"b6",
          4239 => x"81",
          4240 => x"b6",
          4241 => x"81",
          4242 => x"f8",
          4243 => x"74",
          4244 => x"5d",
          4245 => x"5e",
          4246 => x"27",
          4247 => x"73",
          4248 => x"73",
          4249 => x"71",
          4250 => x"5a",
          4251 => x"80",
          4252 => x"38",
          4253 => x"f8",
          4254 => x"0b",
          4255 => x"34",
          4256 => x"33",
          4257 => x"71",
          4258 => x"71",
          4259 => x"71",
          4260 => x"56",
          4261 => x"76",
          4262 => x"ae",
          4263 => x"39",
          4264 => x"38",
          4265 => x"33",
          4266 => x"06",
          4267 => x"11",
          4268 => x"33",
          4269 => x"11",
          4270 => x"80",
          4271 => x"5b",
          4272 => x"86",
          4273 => x"70",
          4274 => x"d8",
          4275 => x"ff",
          4276 => x"d7",
          4277 => x"ff",
          4278 => x"92",
          4279 => x"ff",
          4280 => x"75",
          4281 => x"5e",
          4282 => x"58",
          4283 => x"57",
          4284 => x"8b",
          4285 => x"31",
          4286 => x"29",
          4287 => x"7d",
          4288 => x"74",
          4289 => x"71",
          4290 => x"83",
          4291 => x"62",
          4292 => x"70",
          4293 => x"5f",
          4294 => x"55",
          4295 => x"85",
          4296 => x"29",
          4297 => x"31",
          4298 => x"06",
          4299 => x"fd",
          4300 => x"83",
          4301 => x"fd",
          4302 => x"f2",
          4303 => x"31",
          4304 => x"fe",
          4305 => x"3d",
          4306 => x"80",
          4307 => x"8a",
          4308 => x"73",
          4309 => x"34",
          4310 => x"86",
          4311 => x"55",
          4312 => x"34",
          4313 => x"34",
          4314 => x"98",
          4315 => x"34",
          4316 => x"86",
          4317 => x"54",
          4318 => x"80",
          4319 => x"80",
          4320 => x"52",
          4321 => x"d8",
          4322 => x"87",
          4323 => x"54",
          4324 => x"56",
          4325 => x"f8",
          4326 => x"84",
          4327 => x"72",
          4328 => x"08",
          4329 => x"06",
          4330 => x"51",
          4331 => x"34",
          4332 => x"cc",
          4333 => x"06",
          4334 => x"53",
          4335 => x"81",
          4336 => x"08",
          4337 => x"88",
          4338 => x"75",
          4339 => x"0b",
          4340 => x"34",
          4341 => x"b8",
          4342 => x"3d",
          4343 => x"b6",
          4344 => x"b8",
          4345 => x"f7",
          4346 => x"af",
          4347 => x"84",
          4348 => x"33",
          4349 => x"33",
          4350 => x"81",
          4351 => x"26",
          4352 => x"84",
          4353 => x"83",
          4354 => x"83",
          4355 => x"72",
          4356 => x"86",
          4357 => x"11",
          4358 => x"22",
          4359 => x"59",
          4360 => x"05",
          4361 => x"ff",
          4362 => x"ea",
          4363 => x"58",
          4364 => x"2e",
          4365 => x"83",
          4366 => x"76",
          4367 => x"83",
          4368 => x"83",
          4369 => x"76",
          4370 => x"ff",
          4371 => x"ff",
          4372 => x"55",
          4373 => x"82",
          4374 => x"19",
          4375 => x"f8",
          4376 => x"f8",
          4377 => x"83",
          4378 => x"84",
          4379 => x"5c",
          4380 => x"74",
          4381 => x"38",
          4382 => x"33",
          4383 => x"54",
          4384 => x"72",
          4385 => x"ac",
          4386 => x"b6",
          4387 => x"55",
          4388 => x"33",
          4389 => x"34",
          4390 => x"05",
          4391 => x"70",
          4392 => x"34",
          4393 => x"84",
          4394 => x"27",
          4395 => x"9f",
          4396 => x"38",
          4397 => x"33",
          4398 => x"15",
          4399 => x"0b",
          4400 => x"34",
          4401 => x"81",
          4402 => x"81",
          4403 => x"9f",
          4404 => x"38",
          4405 => x"33",
          4406 => x"75",
          4407 => x"23",
          4408 => x"81",
          4409 => x"83",
          4410 => x"54",
          4411 => x"26",
          4412 => x"72",
          4413 => x"05",
          4414 => x"33",
          4415 => x"58",
          4416 => x"55",
          4417 => x"80",
          4418 => x"b0",
          4419 => x"ff",
          4420 => x"ff",
          4421 => x"29",
          4422 => x"54",
          4423 => x"27",
          4424 => x"97",
          4425 => x"e0",
          4426 => x"53",
          4427 => x"13",
          4428 => x"81",
          4429 => x"73",
          4430 => x"55",
          4431 => x"81",
          4432 => x"81",
          4433 => x"d8",
          4434 => x"d7",
          4435 => x"29",
          4436 => x"5a",
          4437 => x"26",
          4438 => x"53",
          4439 => x"e4",
          4440 => x"0d",
          4441 => x"f8",
          4442 => x"f8",
          4443 => x"83",
          4444 => x"84",
          4445 => x"5c",
          4446 => x"7a",
          4447 => x"38",
          4448 => x"fe",
          4449 => x"81",
          4450 => x"05",
          4451 => x"33",
          4452 => x"75",
          4453 => x"06",
          4454 => x"73",
          4455 => x"05",
          4456 => x"33",
          4457 => x"78",
          4458 => x"56",
          4459 => x"73",
          4460 => x"ae",
          4461 => x"90",
          4462 => x"b6",
          4463 => x"31",
          4464 => x"a0",
          4465 => x"16",
          4466 => x"70",
          4467 => x"34",
          4468 => x"72",
          4469 => x"8a",
          4470 => x"e0",
          4471 => x"75",
          4472 => x"05",
          4473 => x"13",
          4474 => x"38",
          4475 => x"80",
          4476 => x"d8",
          4477 => x"fe",
          4478 => x"f8",
          4479 => x"59",
          4480 => x"19",
          4481 => x"84",
          4482 => x"59",
          4483 => x"fc",
          4484 => x"02",
          4485 => x"05",
          4486 => x"70",
          4487 => x"38",
          4488 => x"83",
          4489 => x"51",
          4490 => x"84",
          4491 => x"51",
          4492 => x"86",
          4493 => x"f8",
          4494 => x"0b",
          4495 => x"0c",
          4496 => x"04",
          4497 => x"f8",
          4498 => x"f8",
          4499 => x"81",
          4500 => x"52",
          4501 => x"e2",
          4502 => x"51",
          4503 => x"94",
          4504 => x"84",
          4505 => x"86",
          4506 => x"83",
          4507 => x"70",
          4508 => x"09",
          4509 => x"72",
          4510 => x"53",
          4511 => x"f8",
          4512 => x"39",
          4513 => x"33",
          4514 => x"b6",
          4515 => x"11",
          4516 => x"70",
          4517 => x"38",
          4518 => x"83",
          4519 => x"80",
          4520 => x"e4",
          4521 => x"0d",
          4522 => x"95",
          4523 => x"31",
          4524 => x"9f",
          4525 => x"54",
          4526 => x"70",
          4527 => x"34",
          4528 => x"b8",
          4529 => x"3d",
          4530 => x"f8",
          4531 => x"05",
          4532 => x"33",
          4533 => x"55",
          4534 => x"25",
          4535 => x"53",
          4536 => x"95",
          4537 => x"84",
          4538 => x"86",
          4539 => x"80",
          4540 => x"95",
          4541 => x"94",
          4542 => x"d7",
          4543 => x"56",
          4544 => x"25",
          4545 => x"81",
          4546 => x"83",
          4547 => x"fe",
          4548 => x"3d",
          4549 => x"05",
          4550 => x"b1",
          4551 => x"70",
          4552 => x"c3",
          4553 => x"70",
          4554 => x"f8",
          4555 => x"80",
          4556 => x"84",
          4557 => x"06",
          4558 => x"2a",
          4559 => x"53",
          4560 => x"f0",
          4561 => x"06",
          4562 => x"f2",
          4563 => x"90",
          4564 => x"84",
          4565 => x"83",
          4566 => x"83",
          4567 => x"81",
          4568 => x"07",
          4569 => x"f8",
          4570 => x"0b",
          4571 => x"0c",
          4572 => x"04",
          4573 => x"33",
          4574 => x"51",
          4575 => x"90",
          4576 => x"83",
          4577 => x"81",
          4578 => x"07",
          4579 => x"f8",
          4580 => x"39",
          4581 => x"83",
          4582 => x"80",
          4583 => x"e4",
          4584 => x"0d",
          4585 => x"90",
          4586 => x"06",
          4587 => x"70",
          4588 => x"34",
          4589 => x"83",
          4590 => x"87",
          4591 => x"83",
          4592 => x"ff",
          4593 => x"f8",
          4594 => x"fd",
          4595 => x"51",
          4596 => x"90",
          4597 => x"39",
          4598 => x"33",
          4599 => x"83",
          4600 => x"83",
          4601 => x"ff",
          4602 => x"f8",
          4603 => x"f9",
          4604 => x"51",
          4605 => x"90",
          4606 => x"39",
          4607 => x"33",
          4608 => x"51",
          4609 => x"90",
          4610 => x"39",
          4611 => x"33",
          4612 => x"80",
          4613 => x"70",
          4614 => x"34",
          4615 => x"83",
          4616 => x"81",
          4617 => x"07",
          4618 => x"f8",
          4619 => x"ba",
          4620 => x"90",
          4621 => x"06",
          4622 => x"51",
          4623 => x"90",
          4624 => x"39",
          4625 => x"33",
          4626 => x"80",
          4627 => x"70",
          4628 => x"34",
          4629 => x"83",
          4630 => x"81",
          4631 => x"07",
          4632 => x"f8",
          4633 => x"82",
          4634 => x"90",
          4635 => x"06",
          4636 => x"f8",
          4637 => x"f2",
          4638 => x"90",
          4639 => x"06",
          4640 => x"70",
          4641 => x"34",
          4642 => x"f3",
          4643 => x"bf",
          4644 => x"84",
          4645 => x"05",
          4646 => x"94",
          4647 => x"93",
          4648 => x"95",
          4649 => x"da",
          4650 => x"5f",
          4651 => x"78",
          4652 => x"a1",
          4653 => x"24",
          4654 => x"81",
          4655 => x"38",
          4656 => x"da",
          4657 => x"84",
          4658 => x"7a",
          4659 => x"34",
          4660 => x"92",
          4661 => x"f8",
          4662 => x"3d",
          4663 => x"83",
          4664 => x"06",
          4665 => x"0b",
          4666 => x"34",
          4667 => x"b6",
          4668 => x"0b",
          4669 => x"34",
          4670 => x"f8",
          4671 => x"0b",
          4672 => x"23",
          4673 => x"b6",
          4674 => x"84",
          4675 => x"56",
          4676 => x"33",
          4677 => x"7c",
          4678 => x"83",
          4679 => x"ff",
          4680 => x"7d",
          4681 => x"34",
          4682 => x"b6",
          4683 => x"83",
          4684 => x"7b",
          4685 => x"23",
          4686 => x"95",
          4687 => x"0d",
          4688 => x"84",
          4689 => x"81",
          4690 => x"dc",
          4691 => x"83",
          4692 => x"a8",
          4693 => x"95",
          4694 => x"83",
          4695 => x"84",
          4696 => x"58",
          4697 => x"33",
          4698 => x"e5",
          4699 => x"55",
          4700 => x"53",
          4701 => x"e2",
          4702 => x"81",
          4703 => x"0b",
          4704 => x"33",
          4705 => x"79",
          4706 => x"79",
          4707 => x"b8",
          4708 => x"53",
          4709 => x"8c",
          4710 => x"ec",
          4711 => x"70",
          4712 => x"84",
          4713 => x"52",
          4714 => x"7a",
          4715 => x"83",
          4716 => x"ff",
          4717 => x"7d",
          4718 => x"34",
          4719 => x"b6",
          4720 => x"83",
          4721 => x"7b",
          4722 => x"23",
          4723 => x"95",
          4724 => x"0d",
          4725 => x"84",
          4726 => x"81",
          4727 => x"dc",
          4728 => x"83",
          4729 => x"a8",
          4730 => x"95",
          4731 => x"83",
          4732 => x"83",
          4733 => x"ff",
          4734 => x"84",
          4735 => x"52",
          4736 => x"51",
          4737 => x"3f",
          4738 => x"f6",
          4739 => x"92",
          4740 => x"84",
          4741 => x"27",
          4742 => x"83",
          4743 => x"33",
          4744 => x"98",
          4745 => x"e0",
          4746 => x"70",
          4747 => x"5a",
          4748 => x"f9",
          4749 => x"02",
          4750 => x"05",
          4751 => x"d8",
          4752 => x"95",
          4753 => x"94",
          4754 => x"29",
          4755 => x"a0",
          4756 => x"f8",
          4757 => x"51",
          4758 => x"7c",
          4759 => x"83",
          4760 => x"83",
          4761 => x"52",
          4762 => x"57",
          4763 => x"2e",
          4764 => x"75",
          4765 => x"f9",
          4766 => x"24",
          4767 => x"75",
          4768 => x"85",
          4769 => x"2e",
          4770 => x"84",
          4771 => x"83",
          4772 => x"83",
          4773 => x"72",
          4774 => x"55",
          4775 => x"b6",
          4776 => x"86",
          4777 => x"14",
          4778 => x"d8",
          4779 => x"95",
          4780 => x"92",
          4781 => x"29",
          4782 => x"56",
          4783 => x"f8",
          4784 => x"83",
          4785 => x"73",
          4786 => x"58",
          4787 => x"90",
          4788 => x"b0",
          4789 => x"84",
          4790 => x"70",
          4791 => x"83",
          4792 => x"83",
          4793 => x"72",
          4794 => x"57",
          4795 => x"57",
          4796 => x"33",
          4797 => x"14",
          4798 => x"70",
          4799 => x"59",
          4800 => x"26",
          4801 => x"84",
          4802 => x"58",
          4803 => x"38",
          4804 => x"72",
          4805 => x"34",
          4806 => x"33",
          4807 => x"2e",
          4808 => x"b6",
          4809 => x"76",
          4810 => x"fb",
          4811 => x"84",
          4812 => x"89",
          4813 => x"75",
          4814 => x"38",
          4815 => x"80",
          4816 => x"8a",
          4817 => x"06",
          4818 => x"81",
          4819 => x"f1",
          4820 => x"0b",
          4821 => x"34",
          4822 => x"83",
          4823 => x"33",
          4824 => x"e0",
          4825 => x"34",
          4826 => x"09",
          4827 => x"89",
          4828 => x"76",
          4829 => x"fd",
          4830 => x"13",
          4831 => x"06",
          4832 => x"83",
          4833 => x"38",
          4834 => x"51",
          4835 => x"81",
          4836 => x"ff",
          4837 => x"83",
          4838 => x"38",
          4839 => x"74",
          4840 => x"34",
          4841 => x"75",
          4842 => x"f9",
          4843 => x"0b",
          4844 => x"0c",
          4845 => x"04",
          4846 => x"2e",
          4847 => x"fd",
          4848 => x"f8",
          4849 => x"81",
          4850 => x"ff",
          4851 => x"83",
          4852 => x"72",
          4853 => x"34",
          4854 => x"51",
          4855 => x"83",
          4856 => x"70",
          4857 => x"55",
          4858 => x"73",
          4859 => x"73",
          4860 => x"f8",
          4861 => x"a0",
          4862 => x"83",
          4863 => x"81",
          4864 => x"ef",
          4865 => x"90",
          4866 => x"75",
          4867 => x"3f",
          4868 => x"e6",
          4869 => x"80",
          4870 => x"84",
          4871 => x"57",
          4872 => x"2e",
          4873 => x"75",
          4874 => x"82",
          4875 => x"2e",
          4876 => x"78",
          4877 => x"d1",
          4878 => x"2e",
          4879 => x"78",
          4880 => x"8f",
          4881 => x"d8",
          4882 => x"94",
          4883 => x"95",
          4884 => x"29",
          4885 => x"5c",
          4886 => x"19",
          4887 => x"a0",
          4888 => x"84",
          4889 => x"83",
          4890 => x"83",
          4891 => x"72",
          4892 => x"5a",
          4893 => x"78",
          4894 => x"18",
          4895 => x"94",
          4896 => x"29",
          4897 => x"5a",
          4898 => x"33",
          4899 => x"b0",
          4900 => x"84",
          4901 => x"70",
          4902 => x"83",
          4903 => x"83",
          4904 => x"72",
          4905 => x"42",
          4906 => x"59",
          4907 => x"33",
          4908 => x"1f",
          4909 => x"70",
          4910 => x"42",
          4911 => x"26",
          4912 => x"84",
          4913 => x"5a",
          4914 => x"38",
          4915 => x"75",
          4916 => x"34",
          4917 => x"b8",
          4918 => x"3d",
          4919 => x"b7",
          4920 => x"38",
          4921 => x"81",
          4922 => x"b8",
          4923 => x"38",
          4924 => x"2e",
          4925 => x"80",
          4926 => x"e0",
          4927 => x"d8",
          4928 => x"94",
          4929 => x"95",
          4930 => x"29",
          4931 => x"40",
          4932 => x"19",
          4933 => x"a0",
          4934 => x"84",
          4935 => x"83",
          4936 => x"83",
          4937 => x"72",
          4938 => x"41",
          4939 => x"78",
          4940 => x"1f",
          4941 => x"94",
          4942 => x"29",
          4943 => x"83",
          4944 => x"86",
          4945 => x"1b",
          4946 => x"d8",
          4947 => x"ff",
          4948 => x"92",
          4949 => x"95",
          4950 => x"29",
          4951 => x"43",
          4952 => x"f8",
          4953 => x"84",
          4954 => x"34",
          4955 => x"77",
          4956 => x"41",
          4957 => x"fe",
          4958 => x"83",
          4959 => x"80",
          4960 => x"e4",
          4961 => x"0d",
          4962 => x"2e",
          4963 => x"78",
          4964 => x"81",
          4965 => x"2e",
          4966 => x"fd",
          4967 => x"0b",
          4968 => x"34",
          4969 => x"b8",
          4970 => x"3d",
          4971 => x"9b",
          4972 => x"38",
          4973 => x"75",
          4974 => x"d0",
          4975 => x"e4",
          4976 => x"59",
          4977 => x"b7",
          4978 => x"84",
          4979 => x"34",
          4980 => x"06",
          4981 => x"84",
          4982 => x"34",
          4983 => x"b8",
          4984 => x"3d",
          4985 => x"9b",
          4986 => x"38",
          4987 => x"b7",
          4988 => x"b6",
          4989 => x"f8",
          4990 => x"f8",
          4991 => x"72",
          4992 => x"40",
          4993 => x"e0",
          4994 => x"a7",
          4995 => x"34",
          4996 => x"33",
          4997 => x"33",
          4998 => x"22",
          4999 => x"12",
          5000 => x"56",
          5001 => x"96",
          5002 => x"f8",
          5003 => x"71",
          5004 => x"57",
          5005 => x"33",
          5006 => x"80",
          5007 => x"b6",
          5008 => x"81",
          5009 => x"f8",
          5010 => x"f8",
          5011 => x"72",
          5012 => x"42",
          5013 => x"83",
          5014 => x"60",
          5015 => x"05",
          5016 => x"58",
          5017 => x"81",
          5018 => x"ea",
          5019 => x"0b",
          5020 => x"34",
          5021 => x"84",
          5022 => x"83",
          5023 => x"70",
          5024 => x"83",
          5025 => x"73",
          5026 => x"86",
          5027 => x"05",
          5028 => x"22",
          5029 => x"72",
          5030 => x"70",
          5031 => x"06",
          5032 => x"33",
          5033 => x"5a",
          5034 => x"2e",
          5035 => x"78",
          5036 => x"ff",
          5037 => x"76",
          5038 => x"76",
          5039 => x"f8",
          5040 => x"90",
          5041 => x"84",
          5042 => x"80",
          5043 => x"e5",
          5044 => x"84",
          5045 => x"80",
          5046 => x"e7",
          5047 => x"84",
          5048 => x"80",
          5049 => x"e4",
          5050 => x"0d",
          5051 => x"94",
          5052 => x"cc",
          5053 => x"95",
          5054 => x"cd",
          5055 => x"93",
          5056 => x"ce",
          5057 => x"84",
          5058 => x"80",
          5059 => x"e4",
          5060 => x"0d",
          5061 => x"ff",
          5062 => x"06",
          5063 => x"83",
          5064 => x"84",
          5065 => x"70",
          5066 => x"83",
          5067 => x"70",
          5068 => x"72",
          5069 => x"86",
          5070 => x"05",
          5071 => x"22",
          5072 => x"7b",
          5073 => x"83",
          5074 => x"83",
          5075 => x"44",
          5076 => x"42",
          5077 => x"81",
          5078 => x"38",
          5079 => x"06",
          5080 => x"56",
          5081 => x"75",
          5082 => x"f8",
          5083 => x"81",
          5084 => x"81",
          5085 => x"81",
          5086 => x"72",
          5087 => x"40",
          5088 => x"80",
          5089 => x"a0",
          5090 => x"84",
          5091 => x"83",
          5092 => x"83",
          5093 => x"72",
          5094 => x"5a",
          5095 => x"a0",
          5096 => x"96",
          5097 => x"f8",
          5098 => x"71",
          5099 => x"5a",
          5100 => x"90",
          5101 => x"b0",
          5102 => x"84",
          5103 => x"70",
          5104 => x"83",
          5105 => x"83",
          5106 => x"72",
          5107 => x"43",
          5108 => x"59",
          5109 => x"33",
          5110 => x"b6",
          5111 => x"1a",
          5112 => x"06",
          5113 => x"7b",
          5114 => x"38",
          5115 => x"33",
          5116 => x"d0",
          5117 => x"58",
          5118 => x"95",
          5119 => x"95",
          5120 => x"ff",
          5121 => x"05",
          5122 => x"39",
          5123 => x"95",
          5124 => x"bd",
          5125 => x"38",
          5126 => x"95",
          5127 => x"b7",
          5128 => x"7e",
          5129 => x"ff",
          5130 => x"75",
          5131 => x"c8",
          5132 => x"10",
          5133 => x"05",
          5134 => x"04",
          5135 => x"f8",
          5136 => x"52",
          5137 => x"9f",
          5138 => x"84",
          5139 => x"9c",
          5140 => x"83",
          5141 => x"84",
          5142 => x"70",
          5143 => x"83",
          5144 => x"70",
          5145 => x"72",
          5146 => x"86",
          5147 => x"05",
          5148 => x"22",
          5149 => x"7b",
          5150 => x"83",
          5151 => x"83",
          5152 => x"46",
          5153 => x"59",
          5154 => x"81",
          5155 => x"38",
          5156 => x"81",
          5157 => x"81",
          5158 => x"81",
          5159 => x"72",
          5160 => x"58",
          5161 => x"80",
          5162 => x"a0",
          5163 => x"84",
          5164 => x"83",
          5165 => x"83",
          5166 => x"72",
          5167 => x"5e",
          5168 => x"a0",
          5169 => x"96",
          5170 => x"f8",
          5171 => x"71",
          5172 => x"5e",
          5173 => x"33",
          5174 => x"80",
          5175 => x"b6",
          5176 => x"81",
          5177 => x"f8",
          5178 => x"f8",
          5179 => x"72",
          5180 => x"44",
          5181 => x"83",
          5182 => x"84",
          5183 => x"34",
          5184 => x"70",
          5185 => x"5b",
          5186 => x"26",
          5187 => x"84",
          5188 => x"58",
          5189 => x"38",
          5190 => x"75",
          5191 => x"34",
          5192 => x"81",
          5193 => x"59",
          5194 => x"f7",
          5195 => x"f8",
          5196 => x"b6",
          5197 => x"f8",
          5198 => x"81",
          5199 => x"81",
          5200 => x"81",
          5201 => x"72",
          5202 => x"5b",
          5203 => x"5b",
          5204 => x"33",
          5205 => x"80",
          5206 => x"b6",
          5207 => x"f8",
          5208 => x"f8",
          5209 => x"71",
          5210 => x"41",
          5211 => x"0b",
          5212 => x"1c",
          5213 => x"94",
          5214 => x"29",
          5215 => x"83",
          5216 => x"86",
          5217 => x"1a",
          5218 => x"d8",
          5219 => x"ff",
          5220 => x"92",
          5221 => x"95",
          5222 => x"29",
          5223 => x"5a",
          5224 => x"f8",
          5225 => x"97",
          5226 => x"60",
          5227 => x"81",
          5228 => x"58",
          5229 => x"fe",
          5230 => x"83",
          5231 => x"fe",
          5232 => x"0b",
          5233 => x"0c",
          5234 => x"b8",
          5235 => x"3d",
          5236 => x"f8",
          5237 => x"59",
          5238 => x"19",
          5239 => x"83",
          5240 => x"70",
          5241 => x"58",
          5242 => x"f9",
          5243 => x"0b",
          5244 => x"34",
          5245 => x"b8",
          5246 => x"3d",
          5247 => x"f8",
          5248 => x"5b",
          5249 => x"1b",
          5250 => x"83",
          5251 => x"84",
          5252 => x"83",
          5253 => x"5b",
          5254 => x"5c",
          5255 => x"84",
          5256 => x"9c",
          5257 => x"53",
          5258 => x"ff",
          5259 => x"84",
          5260 => x"80",
          5261 => x"38",
          5262 => x"33",
          5263 => x"5a",
          5264 => x"e5",
          5265 => x"83",
          5266 => x"02",
          5267 => x"22",
          5268 => x"b8",
          5269 => x"cf",
          5270 => x"96",
          5271 => x"84",
          5272 => x"33",
          5273 => x"f8",
          5274 => x"b6",
          5275 => x"f8",
          5276 => x"5b",
          5277 => x"39",
          5278 => x"33",
          5279 => x"33",
          5280 => x"33",
          5281 => x"05",
          5282 => x"84",
          5283 => x"33",
          5284 => x"a0",
          5285 => x"84",
          5286 => x"83",
          5287 => x"83",
          5288 => x"72",
          5289 => x"5a",
          5290 => x"78",
          5291 => x"18",
          5292 => x"94",
          5293 => x"29",
          5294 => x"83",
          5295 => x"60",
          5296 => x"80",
          5297 => x"b6",
          5298 => x"81",
          5299 => x"f8",
          5300 => x"f8",
          5301 => x"72",
          5302 => x"5f",
          5303 => x"83",
          5304 => x"84",
          5305 => x"34",
          5306 => x"81",
          5307 => x"58",
          5308 => x"90",
          5309 => x"b6",
          5310 => x"77",
          5311 => x"ff",
          5312 => x"83",
          5313 => x"80",
          5314 => x"e0",
          5315 => x"db",
          5316 => x"80",
          5317 => x"38",
          5318 => x"33",
          5319 => x"b4",
          5320 => x"81",
          5321 => x"3f",
          5322 => x"b8",
          5323 => x"3d",
          5324 => x"b8",
          5325 => x"f8",
          5326 => x"b8",
          5327 => x"f8",
          5328 => x"b8",
          5329 => x"76",
          5330 => x"23",
          5331 => x"83",
          5332 => x"84",
          5333 => x"83",
          5334 => x"84",
          5335 => x"83",
          5336 => x"84",
          5337 => x"ff",
          5338 => x"b7",
          5339 => x"7a",
          5340 => x"93",
          5341 => x"b8",
          5342 => x"86",
          5343 => x"06",
          5344 => x"83",
          5345 => x"81",
          5346 => x"f8",
          5347 => x"05",
          5348 => x"83",
          5349 => x"94",
          5350 => x"57",
          5351 => x"3f",
          5352 => x"ff",
          5353 => x"b8",
          5354 => x"ff",
          5355 => x"e8",
          5356 => x"05",
          5357 => x"24",
          5358 => x"76",
          5359 => x"c8",
          5360 => x"ce",
          5361 => x"39",
          5362 => x"b7",
          5363 => x"58",
          5364 => x"06",
          5365 => x"27",
          5366 => x"77",
          5367 => x"b8",
          5368 => x"33",
          5369 => x"b1",
          5370 => x"38",
          5371 => x"83",
          5372 => x"5f",
          5373 => x"84",
          5374 => x"5e",
          5375 => x"8f",
          5376 => x"f8",
          5377 => x"b8",
          5378 => x"71",
          5379 => x"70",
          5380 => x"06",
          5381 => x"5e",
          5382 => x"f8",
          5383 => x"e7",
          5384 => x"e5",
          5385 => x"80",
          5386 => x"38",
          5387 => x"33",
          5388 => x"81",
          5389 => x"b6",
          5390 => x"57",
          5391 => x"27",
          5392 => x"75",
          5393 => x"34",
          5394 => x"80",
          5395 => x"95",
          5396 => x"94",
          5397 => x"ff",
          5398 => x"7b",
          5399 => x"a7",
          5400 => x"56",
          5401 => x"94",
          5402 => x"39",
          5403 => x"f8",
          5404 => x"f8",
          5405 => x"b6",
          5406 => x"05",
          5407 => x"76",
          5408 => x"38",
          5409 => x"75",
          5410 => x"34",
          5411 => x"84",
          5412 => x"40",
          5413 => x"8d",
          5414 => x"f8",
          5415 => x"b8",
          5416 => x"71",
          5417 => x"70",
          5418 => x"06",
          5419 => x"42",
          5420 => x"f8",
          5421 => x"cf",
          5422 => x"e5",
          5423 => x"80",
          5424 => x"38",
          5425 => x"22",
          5426 => x"2e",
          5427 => x"fc",
          5428 => x"b6",
          5429 => x"f8",
          5430 => x"f8",
          5431 => x"71",
          5432 => x"a7",
          5433 => x"83",
          5434 => x"43",
          5435 => x"71",
          5436 => x"70",
          5437 => x"06",
          5438 => x"08",
          5439 => x"80",
          5440 => x"5d",
          5441 => x"82",
          5442 => x"bf",
          5443 => x"83",
          5444 => x"fb",
          5445 => x"b7",
          5446 => x"79",
          5447 => x"e7",
          5448 => x"b8",
          5449 => x"99",
          5450 => x"06",
          5451 => x"81",
          5452 => x"e9",
          5453 => x"39",
          5454 => x"33",
          5455 => x"2e",
          5456 => x"84",
          5457 => x"83",
          5458 => x"5d",
          5459 => x"b6",
          5460 => x"11",
          5461 => x"75",
          5462 => x"38",
          5463 => x"83",
          5464 => x"fb",
          5465 => x"b7",
          5466 => x"76",
          5467 => x"c8",
          5468 => x"b9",
          5469 => x"94",
          5470 => x"05",
          5471 => x"33",
          5472 => x"41",
          5473 => x"25",
          5474 => x"57",
          5475 => x"94",
          5476 => x"39",
          5477 => x"51",
          5478 => x"3f",
          5479 => x"b7",
          5480 => x"57",
          5481 => x"8b",
          5482 => x"10",
          5483 => x"05",
          5484 => x"5a",
          5485 => x"51",
          5486 => x"3f",
          5487 => x"81",
          5488 => x"b7",
          5489 => x"58",
          5490 => x"82",
          5491 => x"e5",
          5492 => x"7d",
          5493 => x"38",
          5494 => x"22",
          5495 => x"26",
          5496 => x"57",
          5497 => x"81",
          5498 => x"d5",
          5499 => x"97",
          5500 => x"e5",
          5501 => x"77",
          5502 => x"38",
          5503 => x"33",
          5504 => x"81",
          5505 => x"b8",
          5506 => x"05",
          5507 => x"06",
          5508 => x"33",
          5509 => x"06",
          5510 => x"43",
          5511 => x"5c",
          5512 => x"27",
          5513 => x"5a",
          5514 => x"92",
          5515 => x"ff",
          5516 => x"58",
          5517 => x"27",
          5518 => x"57",
          5519 => x"94",
          5520 => x"d8",
          5521 => x"57",
          5522 => x"27",
          5523 => x"7a",
          5524 => x"f8",
          5525 => x"af",
          5526 => x"e5",
          5527 => x"80",
          5528 => x"38",
          5529 => x"33",
          5530 => x"33",
          5531 => x"7f",
          5532 => x"38",
          5533 => x"33",
          5534 => x"33",
          5535 => x"06",
          5536 => x"33",
          5537 => x"11",
          5538 => x"80",
          5539 => x"92",
          5540 => x"71",
          5541 => x"70",
          5542 => x"06",
          5543 => x"33",
          5544 => x"59",
          5545 => x"81",
          5546 => x"38",
          5547 => x"ff",
          5548 => x"31",
          5549 => x"7c",
          5550 => x"38",
          5551 => x"33",
          5552 => x"27",
          5553 => x"ff",
          5554 => x"83",
          5555 => x"7c",
          5556 => x"70",
          5557 => x"57",
          5558 => x"8e",
          5559 => x"b6",
          5560 => x"76",
          5561 => x"ee",
          5562 => x"56",
          5563 => x"94",
          5564 => x"ff",
          5565 => x"92",
          5566 => x"80",
          5567 => x"26",
          5568 => x"77",
          5569 => x"7e",
          5570 => x"71",
          5571 => x"5e",
          5572 => x"86",
          5573 => x"5b",
          5574 => x"80",
          5575 => x"06",
          5576 => x"06",
          5577 => x"1d",
          5578 => x"5c",
          5579 => x"f7",
          5580 => x"97",
          5581 => x"e0",
          5582 => x"5f",
          5583 => x"1f",
          5584 => x"81",
          5585 => x"76",
          5586 => x"58",
          5587 => x"81",
          5588 => x"81",
          5589 => x"d8",
          5590 => x"d7",
          5591 => x"29",
          5592 => x"5e",
          5593 => x"27",
          5594 => x"e0",
          5595 => x"5f",
          5596 => x"1f",
          5597 => x"81",
          5598 => x"76",
          5599 => x"58",
          5600 => x"81",
          5601 => x"81",
          5602 => x"d8",
          5603 => x"d7",
          5604 => x"29",
          5605 => x"5e",
          5606 => x"26",
          5607 => x"f6",
          5608 => x"b7",
          5609 => x"75",
          5610 => x"e0",
          5611 => x"84",
          5612 => x"51",
          5613 => x"f6",
          5614 => x"0b",
          5615 => x"33",
          5616 => x"b7",
          5617 => x"59",
          5618 => x"78",
          5619 => x"84",
          5620 => x"56",
          5621 => x"09",
          5622 => x"be",
          5623 => x"95",
          5624 => x"81",
          5625 => x"f8",
          5626 => x"43",
          5627 => x"ff",
          5628 => x"38",
          5629 => x"33",
          5630 => x"26",
          5631 => x"7e",
          5632 => x"56",
          5633 => x"f5",
          5634 => x"76",
          5635 => x"27",
          5636 => x"f5",
          5637 => x"10",
          5638 => x"90",
          5639 => x"86",
          5640 => x"11",
          5641 => x"5a",
          5642 => x"80",
          5643 => x"06",
          5644 => x"75",
          5645 => x"79",
          5646 => x"76",
          5647 => x"83",
          5648 => x"70",
          5649 => x"90",
          5650 => x"88",
          5651 => x"07",
          5652 => x"52",
          5653 => x"7a",
          5654 => x"80",
          5655 => x"05",
          5656 => x"76",
          5657 => x"58",
          5658 => x"26",
          5659 => x"b6",
          5660 => x"b6",
          5661 => x"5f",
          5662 => x"06",
          5663 => x"06",
          5664 => x"22",
          5665 => x"64",
          5666 => x"59",
          5667 => x"26",
          5668 => x"78",
          5669 => x"7b",
          5670 => x"57",
          5671 => x"1d",
          5672 => x"76",
          5673 => x"38",
          5674 => x"33",
          5675 => x"18",
          5676 => x"0b",
          5677 => x"34",
          5678 => x"81",
          5679 => x"81",
          5680 => x"76",
          5681 => x"38",
          5682 => x"e0",
          5683 => x"78",
          5684 => x"5a",
          5685 => x"57",
          5686 => x"d6",
          5687 => x"39",
          5688 => x"81",
          5689 => x"58",
          5690 => x"83",
          5691 => x"70",
          5692 => x"71",
          5693 => x"f0",
          5694 => x"2a",
          5695 => x"57",
          5696 => x"2e",
          5697 => x"be",
          5698 => x"0b",
          5699 => x"34",
          5700 => x"81",
          5701 => x"56",
          5702 => x"83",
          5703 => x"33",
          5704 => x"e0",
          5705 => x"34",
          5706 => x"33",
          5707 => x"33",
          5708 => x"22",
          5709 => x"33",
          5710 => x"5d",
          5711 => x"83",
          5712 => x"87",
          5713 => x"83",
          5714 => x"81",
          5715 => x"ff",
          5716 => x"f4",
          5717 => x"f8",
          5718 => x"fd",
          5719 => x"56",
          5720 => x"90",
          5721 => x"83",
          5722 => x"81",
          5723 => x"07",
          5724 => x"f8",
          5725 => x"39",
          5726 => x"33",
          5727 => x"81",
          5728 => x"83",
          5729 => x"c3",
          5730 => x"90",
          5731 => x"06",
          5732 => x"75",
          5733 => x"34",
          5734 => x"80",
          5735 => x"f8",
          5736 => x"18",
          5737 => x"06",
          5738 => x"a4",
          5739 => x"90",
          5740 => x"06",
          5741 => x"f8",
          5742 => x"8f",
          5743 => x"90",
          5744 => x"06",
          5745 => x"75",
          5746 => x"34",
          5747 => x"83",
          5748 => x"81",
          5749 => x"e0",
          5750 => x"83",
          5751 => x"fe",
          5752 => x"f8",
          5753 => x"cf",
          5754 => x"07",
          5755 => x"f8",
          5756 => x"d7",
          5757 => x"90",
          5758 => x"06",
          5759 => x"75",
          5760 => x"34",
          5761 => x"83",
          5762 => x"81",
          5763 => x"07",
          5764 => x"f8",
          5765 => x"b3",
          5766 => x"90",
          5767 => x"06",
          5768 => x"75",
          5769 => x"34",
          5770 => x"83",
          5771 => x"81",
          5772 => x"07",
          5773 => x"f8",
          5774 => x"8f",
          5775 => x"90",
          5776 => x"06",
          5777 => x"f8",
          5778 => x"ff",
          5779 => x"90",
          5780 => x"07",
          5781 => x"f8",
          5782 => x"ef",
          5783 => x"90",
          5784 => x"07",
          5785 => x"f8",
          5786 => x"df",
          5787 => x"90",
          5788 => x"06",
          5789 => x"56",
          5790 => x"90",
          5791 => x"39",
          5792 => x"33",
          5793 => x"b0",
          5794 => x"83",
          5795 => x"fd",
          5796 => x"0b",
          5797 => x"34",
          5798 => x"51",
          5799 => x"ec",
          5800 => x"b8",
          5801 => x"f8",
          5802 => x"b8",
          5803 => x"f8",
          5804 => x"b8",
          5805 => x"78",
          5806 => x"23",
          5807 => x"b7",
          5808 => x"c7",
          5809 => x"84",
          5810 => x"80",
          5811 => x"e4",
          5812 => x"0d",
          5813 => x"f8",
          5814 => x"f8",
          5815 => x"81",
          5816 => x"ff",
          5817 => x"cf",
          5818 => x"e8",
          5819 => x"dc",
          5820 => x"05",
          5821 => x"8e",
          5822 => x"e4",
          5823 => x"84",
          5824 => x"84",
          5825 => x"80",
          5826 => x"e4",
          5827 => x"84",
          5828 => x"9c",
          5829 => x"77",
          5830 => x"34",
          5831 => x"84",
          5832 => x"81",
          5833 => x"7a",
          5834 => x"34",
          5835 => x"fe",
          5836 => x"80",
          5837 => x"84",
          5838 => x"23",
          5839 => x"b7",
          5840 => x"39",
          5841 => x"f8",
          5842 => x"52",
          5843 => x"97",
          5844 => x"95",
          5845 => x"ff",
          5846 => x"05",
          5847 => x"39",
          5848 => x"f8",
          5849 => x"52",
          5850 => x"fb",
          5851 => x"39",
          5852 => x"eb",
          5853 => x"8f",
          5854 => x"95",
          5855 => x"70",
          5856 => x"2c",
          5857 => x"5f",
          5858 => x"39",
          5859 => x"51",
          5860 => x"b6",
          5861 => x"75",
          5862 => x"eb",
          5863 => x"f8",
          5864 => x"e3",
          5865 => x"94",
          5866 => x"70",
          5867 => x"2c",
          5868 => x"40",
          5869 => x"39",
          5870 => x"33",
          5871 => x"b6",
          5872 => x"11",
          5873 => x"75",
          5874 => x"c0",
          5875 => x"f3",
          5876 => x"b6",
          5877 => x"81",
          5878 => x"5c",
          5879 => x"ee",
          5880 => x"f8",
          5881 => x"b6",
          5882 => x"81",
          5883 => x"f8",
          5884 => x"74",
          5885 => x"a7",
          5886 => x"83",
          5887 => x"5f",
          5888 => x"29",
          5889 => x"ff",
          5890 => x"f6",
          5891 => x"5b",
          5892 => x"5d",
          5893 => x"81",
          5894 => x"83",
          5895 => x"ff",
          5896 => x"80",
          5897 => x"89",
          5898 => x"d7",
          5899 => x"76",
          5900 => x"38",
          5901 => x"75",
          5902 => x"23",
          5903 => x"06",
          5904 => x"57",
          5905 => x"83",
          5906 => x"b6",
          5907 => x"76",
          5908 => x"ec",
          5909 => x"56",
          5910 => x"94",
          5911 => x"ff",
          5912 => x"92",
          5913 => x"80",
          5914 => x"26",
          5915 => x"77",
          5916 => x"7e",
          5917 => x"71",
          5918 => x"5e",
          5919 => x"86",
          5920 => x"5b",
          5921 => x"80",
          5922 => x"06",
          5923 => x"06",
          5924 => x"1d",
          5925 => x"5d",
          5926 => x"ec",
          5927 => x"97",
          5928 => x"e0",
          5929 => x"5e",
          5930 => x"1e",
          5931 => x"81",
          5932 => x"76",
          5933 => x"58",
          5934 => x"81",
          5935 => x"81",
          5936 => x"d8",
          5937 => x"d7",
          5938 => x"29",
          5939 => x"5d",
          5940 => x"27",
          5941 => x"e0",
          5942 => x"5e",
          5943 => x"1e",
          5944 => x"81",
          5945 => x"76",
          5946 => x"58",
          5947 => x"81",
          5948 => x"81",
          5949 => x"d8",
          5950 => x"d7",
          5951 => x"29",
          5952 => x"5d",
          5953 => x"26",
          5954 => x"eb",
          5955 => x"f8",
          5956 => x"5c",
          5957 => x"1c",
          5958 => x"83",
          5959 => x"84",
          5960 => x"83",
          5961 => x"84",
          5962 => x"5f",
          5963 => x"fd",
          5964 => x"eb",
          5965 => x"b6",
          5966 => x"81",
          5967 => x"11",
          5968 => x"76",
          5969 => x"38",
          5970 => x"83",
          5971 => x"77",
          5972 => x"ff",
          5973 => x"80",
          5974 => x"38",
          5975 => x"83",
          5976 => x"84",
          5977 => x"70",
          5978 => x"ff",
          5979 => x"56",
          5980 => x"eb",
          5981 => x"56",
          5982 => x"95",
          5983 => x"39",
          5984 => x"33",
          5985 => x"b6",
          5986 => x"11",
          5987 => x"75",
          5988 => x"ca",
          5989 => x"ef",
          5990 => x"81",
          5991 => x"06",
          5992 => x"83",
          5993 => x"70",
          5994 => x"83",
          5995 => x"7a",
          5996 => x"57",
          5997 => x"09",
          5998 => x"b8",
          5999 => x"39",
          6000 => x"75",
          6001 => x"34",
          6002 => x"ff",
          6003 => x"83",
          6004 => x"fc",
          6005 => x"7b",
          6006 => x"83",
          6007 => x"f2",
          6008 => x"7d",
          6009 => x"7a",
          6010 => x"38",
          6011 => x"81",
          6012 => x"83",
          6013 => x"77",
          6014 => x"59",
          6015 => x"26",
          6016 => x"80",
          6017 => x"05",
          6018 => x"f8",
          6019 => x"70",
          6020 => x"34",
          6021 => x"d4",
          6022 => x"39",
          6023 => x"56",
          6024 => x"92",
          6025 => x"39",
          6026 => x"f8",
          6027 => x"ad",
          6028 => x"f8",
          6029 => x"84",
          6030 => x"83",
          6031 => x"f1",
          6032 => x"0b",
          6033 => x"34",
          6034 => x"83",
          6035 => x"33",
          6036 => x"e0",
          6037 => x"34",
          6038 => x"f6",
          6039 => x"a7",
          6040 => x"0d",
          6041 => x"33",
          6042 => x"33",
          6043 => x"80",
          6044 => x"73",
          6045 => x"3f",
          6046 => x"b8",
          6047 => x"3d",
          6048 => x"52",
          6049 => x"ab",
          6050 => x"84",
          6051 => x"85",
          6052 => x"f3",
          6053 => x"bf",
          6054 => x"ff",
          6055 => x"e8",
          6056 => x"ff",
          6057 => x"c8",
          6058 => x"55",
          6059 => x"80",
          6060 => x"38",
          6061 => x"75",
          6062 => x"34",
          6063 => x"84",
          6064 => x"8f",
          6065 => x"83",
          6066 => x"54",
          6067 => x"80",
          6068 => x"73",
          6069 => x"30",
          6070 => x"09",
          6071 => x"56",
          6072 => x"72",
          6073 => x"0c",
          6074 => x"54",
          6075 => x"09",
          6076 => x"38",
          6077 => x"83",
          6078 => x"70",
          6079 => x"07",
          6080 => x"79",
          6081 => x"c4",
          6082 => x"d8",
          6083 => x"95",
          6084 => x"94",
          6085 => x"29",
          6086 => x"a0",
          6087 => x"f8",
          6088 => x"59",
          6089 => x"29",
          6090 => x"ff",
          6091 => x"f6",
          6092 => x"59",
          6093 => x"81",
          6094 => x"38",
          6095 => x"73",
          6096 => x"80",
          6097 => x"87",
          6098 => x"0c",
          6099 => x"88",
          6100 => x"80",
          6101 => x"86",
          6102 => x"08",
          6103 => x"f4",
          6104 => x"81",
          6105 => x"ff",
          6106 => x"81",
          6107 => x"cf",
          6108 => x"83",
          6109 => x"33",
          6110 => x"06",
          6111 => x"16",
          6112 => x"55",
          6113 => x"85",
          6114 => x"81",
          6115 => x"b4",
          6116 => x"f6",
          6117 => x"75",
          6118 => x"5a",
          6119 => x"2e",
          6120 => x"75",
          6121 => x"15",
          6122 => x"84",
          6123 => x"f6",
          6124 => x"81",
          6125 => x"ff",
          6126 => x"89",
          6127 => x"b3",
          6128 => x"8c",
          6129 => x"2b",
          6130 => x"58",
          6131 => x"83",
          6132 => x"73",
          6133 => x"70",
          6134 => x"32",
          6135 => x"51",
          6136 => x"80",
          6137 => x"38",
          6138 => x"f6",
          6139 => x"09",
          6140 => x"72",
          6141 => x"e4",
          6142 => x"83",
          6143 => x"80",
          6144 => x"bd",
          6145 => x"c4",
          6146 => x"be",
          6147 => x"f6",
          6148 => x"f6",
          6149 => x"5d",
          6150 => x"5e",
          6151 => x"98",
          6152 => x"74",
          6153 => x"8d",
          6154 => x"ac",
          6155 => x"73",
          6156 => x"82",
          6157 => x"a2",
          6158 => x"72",
          6159 => x"8b",
          6160 => x"ac",
          6161 => x"73",
          6162 => x"74",
          6163 => x"54",
          6164 => x"2e",
          6165 => x"f6",
          6166 => x"53",
          6167 => x"81",
          6168 => x"81",
          6169 => x"72",
          6170 => x"84",
          6171 => x"f6",
          6172 => x"54",
          6173 => x"84",
          6174 => x"f6",
          6175 => x"e8",
          6176 => x"98",
          6177 => x"54",
          6178 => x"83",
          6179 => x"0b",
          6180 => x"9c",
          6181 => x"b8",
          6182 => x"16",
          6183 => x"06",
          6184 => x"76",
          6185 => x"38",
          6186 => x"bf",
          6187 => x"f6",
          6188 => x"9e",
          6189 => x"9c",
          6190 => x"38",
          6191 => x"83",
          6192 => x"5a",
          6193 => x"83",
          6194 => x"54",
          6195 => x"91",
          6196 => x"14",
          6197 => x"9c",
          6198 => x"7d",
          6199 => x"dc",
          6200 => x"83",
          6201 => x"54",
          6202 => x"2e",
          6203 => x"54",
          6204 => x"ea",
          6205 => x"98",
          6206 => x"f6",
          6207 => x"81",
          6208 => x"77",
          6209 => x"38",
          6210 => x"17",
          6211 => x"b6",
          6212 => x"76",
          6213 => x"54",
          6214 => x"83",
          6215 => x"53",
          6216 => x"82",
          6217 => x"81",
          6218 => x"38",
          6219 => x"34",
          6220 => x"fc",
          6221 => x"58",
          6222 => x"80",
          6223 => x"83",
          6224 => x"2e",
          6225 => x"77",
          6226 => x"06",
          6227 => x"7d",
          6228 => x"ed",
          6229 => x"2e",
          6230 => x"79",
          6231 => x"59",
          6232 => x"75",
          6233 => x"54",
          6234 => x"a1",
          6235 => x"2e",
          6236 => x"17",
          6237 => x"06",
          6238 => x"fe",
          6239 => x"27",
          6240 => x"57",
          6241 => x"54",
          6242 => x"e1",
          6243 => x"10",
          6244 => x"05",
          6245 => x"2b",
          6246 => x"f2",
          6247 => x"33",
          6248 => x"78",
          6249 => x"9c",
          6250 => x"b8",
          6251 => x"ea",
          6252 => x"7d",
          6253 => x"a8",
          6254 => x"ff",
          6255 => x"a0",
          6256 => x"ff",
          6257 => x"ff",
          6258 => x"38",
          6259 => x"b6",
          6260 => x"54",
          6261 => x"83",
          6262 => x"82",
          6263 => x"70",
          6264 => x"07",
          6265 => x"7d",
          6266 => x"83",
          6267 => x"06",
          6268 => x"78",
          6269 => x"c6",
          6270 => x"72",
          6271 => x"83",
          6272 => x"70",
          6273 => x"78",
          6274 => x"ba",
          6275 => x"70",
          6276 => x"54",
          6277 => x"27",
          6278 => x"b6",
          6279 => x"72",
          6280 => x"9a",
          6281 => x"dc",
          6282 => x"f9",
          6283 => x"81",
          6284 => x"82",
          6285 => x"3f",
          6286 => x"e4",
          6287 => x"0d",
          6288 => x"34",
          6289 => x"f9",
          6290 => x"81",
          6291 => x"38",
          6292 => x"14",
          6293 => x"5b",
          6294 => x"ac",
          6295 => x"c9",
          6296 => x"83",
          6297 => x"34",
          6298 => x"f6",
          6299 => x"ff",
          6300 => x"a2",
          6301 => x"b1",
          6302 => x"ff",
          6303 => x"81",
          6304 => x"96",
          6305 => x"ac",
          6306 => x"81",
          6307 => x"8a",
          6308 => x"ff",
          6309 => x"81",
          6310 => x"06",
          6311 => x"83",
          6312 => x"81",
          6313 => x"c0",
          6314 => x"54",
          6315 => x"27",
          6316 => x"87",
          6317 => x"08",
          6318 => x"0c",
          6319 => x"06",
          6320 => x"39",
          6321 => x"f6",
          6322 => x"f9",
          6323 => x"83",
          6324 => x"73",
          6325 => x"53",
          6326 => x"38",
          6327 => x"be",
          6328 => x"83",
          6329 => x"83",
          6330 => x"83",
          6331 => x"70",
          6332 => x"33",
          6333 => x"33",
          6334 => x"5e",
          6335 => x"fa",
          6336 => x"82",
          6337 => x"06",
          6338 => x"7a",
          6339 => x"2e",
          6340 => x"79",
          6341 => x"81",
          6342 => x"38",
          6343 => x"ef",
          6344 => x"f0",
          6345 => x"39",
          6346 => x"b6",
          6347 => x"54",
          6348 => x"81",
          6349 => x"b6",
          6350 => x"59",
          6351 => x"80",
          6352 => x"da",
          6353 => x"76",
          6354 => x"54",
          6355 => x"da",
          6356 => x"f7",
          6357 => x"53",
          6358 => x"08",
          6359 => x"83",
          6360 => x"83",
          6361 => x"f6",
          6362 => x"b6",
          6363 => x"81",
          6364 => x"11",
          6365 => x"80",
          6366 => x"38",
          6367 => x"83",
          6368 => x"73",
          6369 => x"ff",
          6370 => x"80",
          6371 => x"38",
          6372 => x"83",
          6373 => x"84",
          6374 => x"70",
          6375 => x"56",
          6376 => x"80",
          6377 => x"38",
          6378 => x"83",
          6379 => x"ff",
          6380 => x"39",
          6381 => x"51",
          6382 => x"3f",
          6383 => x"aa",
          6384 => x"fc",
          6385 => x"14",
          6386 => x"f6",
          6387 => x"de",
          6388 => x"0b",
          6389 => x"34",
          6390 => x"33",
          6391 => x"39",
          6392 => x"81",
          6393 => x"3f",
          6394 => x"04",
          6395 => x"80",
          6396 => x"f0",
          6397 => x"02",
          6398 => x"82",
          6399 => x"f2",
          6400 => x"80",
          6401 => x"85",
          6402 => x"f0",
          6403 => x"fe",
          6404 => x"34",
          6405 => x"f0",
          6406 => x"87",
          6407 => x"08",
          6408 => x"08",
          6409 => x"90",
          6410 => x"c0",
          6411 => x"52",
          6412 => x"9c",
          6413 => x"72",
          6414 => x"81",
          6415 => x"c0",
          6416 => x"56",
          6417 => x"27",
          6418 => x"81",
          6419 => x"38",
          6420 => x"a4",
          6421 => x"55",
          6422 => x"80",
          6423 => x"55",
          6424 => x"80",
          6425 => x"c0",
          6426 => x"80",
          6427 => x"53",
          6428 => x"9c",
          6429 => x"c0",
          6430 => x"55",
          6431 => x"f6",
          6432 => x"33",
          6433 => x"9c",
          6434 => x"70",
          6435 => x"38",
          6436 => x"2e",
          6437 => x"c0",
          6438 => x"55",
          6439 => x"83",
          6440 => x"71",
          6441 => x"70",
          6442 => x"57",
          6443 => x"2e",
          6444 => x"81",
          6445 => x"71",
          6446 => x"74",
          6447 => x"38",
          6448 => x"e4",
          6449 => x"0d",
          6450 => x"84",
          6451 => x"88",
          6452 => x"fa",
          6453 => x"02",
          6454 => x"05",
          6455 => x"80",
          6456 => x"f0",
          6457 => x"2b",
          6458 => x"80",
          6459 => x"98",
          6460 => x"55",
          6461 => x"83",
          6462 => x"90",
          6463 => x"84",
          6464 => x"90",
          6465 => x"85",
          6466 => x"86",
          6467 => x"f2",
          6468 => x"74",
          6469 => x"83",
          6470 => x"51",
          6471 => x"34",
          6472 => x"f2",
          6473 => x"56",
          6474 => x"15",
          6475 => x"86",
          6476 => x"34",
          6477 => x"9c",
          6478 => x"f0",
          6479 => x"ce",
          6480 => x"87",
          6481 => x"08",
          6482 => x"98",
          6483 => x"70",
          6484 => x"38",
          6485 => x"87",
          6486 => x"08",
          6487 => x"73",
          6488 => x"71",
          6489 => x"db",
          6490 => x"98",
          6491 => x"ff",
          6492 => x"27",
          6493 => x"71",
          6494 => x"2e",
          6495 => x"87",
          6496 => x"08",
          6497 => x"05",
          6498 => x"98",
          6499 => x"87",
          6500 => x"08",
          6501 => x"2e",
          6502 => x"14",
          6503 => x"98",
          6504 => x"52",
          6505 => x"87",
          6506 => x"ff",
          6507 => x"87",
          6508 => x"08",
          6509 => x"26",
          6510 => x"52",
          6511 => x"16",
          6512 => x"06",
          6513 => x"80",
          6514 => x"38",
          6515 => x"06",
          6516 => x"d4",
          6517 => x"70",
          6518 => x"56",
          6519 => x"80",
          6520 => x"84",
          6521 => x"52",
          6522 => x"27",
          6523 => x"70",
          6524 => x"33",
          6525 => x"05",
          6526 => x"71",
          6527 => x"76",
          6528 => x"0c",
          6529 => x"04",
          6530 => x"b8",
          6531 => x"3d",
          6532 => x"51",
          6533 => x"3d",
          6534 => x"84",
          6535 => x"33",
          6536 => x"0b",
          6537 => x"08",
          6538 => x"87",
          6539 => x"06",
          6540 => x"2a",
          6541 => x"55",
          6542 => x"15",
          6543 => x"2a",
          6544 => x"15",
          6545 => x"2a",
          6546 => x"15",
          6547 => x"15",
          6548 => x"f2",
          6549 => x"c6",
          6550 => x"13",
          6551 => x"51",
          6552 => x"97",
          6553 => x"81",
          6554 => x"72",
          6555 => x"54",
          6556 => x"26",
          6557 => x"f2",
          6558 => x"74",
          6559 => x"83",
          6560 => x"55",
          6561 => x"34",
          6562 => x"f2",
          6563 => x"56",
          6564 => x"15",
          6565 => x"86",
          6566 => x"34",
          6567 => x"9c",
          6568 => x"f0",
          6569 => x"ce",
          6570 => x"87",
          6571 => x"08",
          6572 => x"98",
          6573 => x"70",
          6574 => x"38",
          6575 => x"87",
          6576 => x"08",
          6577 => x"73",
          6578 => x"71",
          6579 => x"db",
          6580 => x"98",
          6581 => x"ff",
          6582 => x"27",
          6583 => x"71",
          6584 => x"2e",
          6585 => x"87",
          6586 => x"08",
          6587 => x"05",
          6588 => x"98",
          6589 => x"87",
          6590 => x"08",
          6591 => x"2e",
          6592 => x"14",
          6593 => x"98",
          6594 => x"52",
          6595 => x"87",
          6596 => x"ff",
          6597 => x"87",
          6598 => x"08",
          6599 => x"26",
          6600 => x"52",
          6601 => x"16",
          6602 => x"06",
          6603 => x"80",
          6604 => x"74",
          6605 => x"52",
          6606 => x"38",
          6607 => x"81",
          6608 => x"73",
          6609 => x"38",
          6610 => x"84",
          6611 => x"88",
          6612 => x"ff",
          6613 => x"fb",
          6614 => x"f2",
          6615 => x"80",
          6616 => x"85",
          6617 => x"f0",
          6618 => x"fe",
          6619 => x"34",
          6620 => x"f0",
          6621 => x"87",
          6622 => x"08",
          6623 => x"08",
          6624 => x"90",
          6625 => x"c0",
          6626 => x"52",
          6627 => x"9c",
          6628 => x"72",
          6629 => x"81",
          6630 => x"c0",
          6631 => x"52",
          6632 => x"27",
          6633 => x"81",
          6634 => x"38",
          6635 => x"a4",
          6636 => x"53",
          6637 => x"80",
          6638 => x"53",
          6639 => x"80",
          6640 => x"c0",
          6641 => x"80",
          6642 => x"53",
          6643 => x"9c",
          6644 => x"c0",
          6645 => x"51",
          6646 => x"f6",
          6647 => x"33",
          6648 => x"9c",
          6649 => x"73",
          6650 => x"38",
          6651 => x"2e",
          6652 => x"c0",
          6653 => x"51",
          6654 => x"83",
          6655 => x"71",
          6656 => x"70",
          6657 => x"57",
          6658 => x"2e",
          6659 => x"81",
          6660 => x"73",
          6661 => x"ff",
          6662 => x"0d",
          6663 => x"51",
          6664 => x"3f",
          6665 => x"04",
          6666 => x"84",
          6667 => x"7a",
          6668 => x"2a",
          6669 => x"ff",
          6670 => x"2b",
          6671 => x"33",
          6672 => x"71",
          6673 => x"83",
          6674 => x"11",
          6675 => x"12",
          6676 => x"2b",
          6677 => x"07",
          6678 => x"53",
          6679 => x"59",
          6680 => x"53",
          6681 => x"81",
          6682 => x"16",
          6683 => x"83",
          6684 => x"8b",
          6685 => x"2b",
          6686 => x"70",
          6687 => x"33",
          6688 => x"71",
          6689 => x"57",
          6690 => x"59",
          6691 => x"71",
          6692 => x"38",
          6693 => x"85",
          6694 => x"8b",
          6695 => x"2b",
          6696 => x"76",
          6697 => x"54",
          6698 => x"86",
          6699 => x"81",
          6700 => x"73",
          6701 => x"84",
          6702 => x"70",
          6703 => x"33",
          6704 => x"71",
          6705 => x"70",
          6706 => x"55",
          6707 => x"77",
          6708 => x"71",
          6709 => x"84",
          6710 => x"16",
          6711 => x"86",
          6712 => x"0b",
          6713 => x"84",
          6714 => x"53",
          6715 => x"34",
          6716 => x"34",
          6717 => x"08",
          6718 => x"81",
          6719 => x"88",
          6720 => x"80",
          6721 => x"88",
          6722 => x"52",
          6723 => x"34",
          6724 => x"34",
          6725 => x"04",
          6726 => x"87",
          6727 => x"8b",
          6728 => x"2b",
          6729 => x"84",
          6730 => x"17",
          6731 => x"2b",
          6732 => x"2a",
          6733 => x"51",
          6734 => x"71",
          6735 => x"72",
          6736 => x"84",
          6737 => x"70",
          6738 => x"33",
          6739 => x"71",
          6740 => x"83",
          6741 => x"5a",
          6742 => x"05",
          6743 => x"87",
          6744 => x"88",
          6745 => x"88",
          6746 => x"59",
          6747 => x"13",
          6748 => x"13",
          6749 => x"d4",
          6750 => x"33",
          6751 => x"71",
          6752 => x"81",
          6753 => x"70",
          6754 => x"5a",
          6755 => x"72",
          6756 => x"13",
          6757 => x"d4",
          6758 => x"70",
          6759 => x"33",
          6760 => x"71",
          6761 => x"74",
          6762 => x"81",
          6763 => x"88",
          6764 => x"83",
          6765 => x"f8",
          6766 => x"7b",
          6767 => x"52",
          6768 => x"5a",
          6769 => x"77",
          6770 => x"73",
          6771 => x"84",
          6772 => x"70",
          6773 => x"81",
          6774 => x"8b",
          6775 => x"2b",
          6776 => x"70",
          6777 => x"33",
          6778 => x"07",
          6779 => x"06",
          6780 => x"5f",
          6781 => x"5a",
          6782 => x"77",
          6783 => x"81",
          6784 => x"b8",
          6785 => x"17",
          6786 => x"83",
          6787 => x"8b",
          6788 => x"2b",
          6789 => x"70",
          6790 => x"33",
          6791 => x"71",
          6792 => x"58",
          6793 => x"5a",
          6794 => x"70",
          6795 => x"e4",
          6796 => x"81",
          6797 => x"88",
          6798 => x"80",
          6799 => x"88",
          6800 => x"54",
          6801 => x"77",
          6802 => x"84",
          6803 => x"70",
          6804 => x"81",
          6805 => x"8b",
          6806 => x"2b",
          6807 => x"82",
          6808 => x"15",
          6809 => x"2b",
          6810 => x"2a",
          6811 => x"52",
          6812 => x"53",
          6813 => x"34",
          6814 => x"34",
          6815 => x"04",
          6816 => x"79",
          6817 => x"08",
          6818 => x"80",
          6819 => x"77",
          6820 => x"38",
          6821 => x"90",
          6822 => x"0d",
          6823 => x"f4",
          6824 => x"d4",
          6825 => x"0b",
          6826 => x"23",
          6827 => x"53",
          6828 => x"ff",
          6829 => x"d3",
          6830 => x"b8",
          6831 => x"76",
          6832 => x"0b",
          6833 => x"84",
          6834 => x"54",
          6835 => x"34",
          6836 => x"15",
          6837 => x"d4",
          6838 => x"86",
          6839 => x"0b",
          6840 => x"84",
          6841 => x"84",
          6842 => x"ff",
          6843 => x"80",
          6844 => x"ff",
          6845 => x"88",
          6846 => x"55",
          6847 => x"17",
          6848 => x"17",
          6849 => x"d0",
          6850 => x"10",
          6851 => x"d4",
          6852 => x"05",
          6853 => x"82",
          6854 => x"0b",
          6855 => x"fe",
          6856 => x"3d",
          6857 => x"80",
          6858 => x"84",
          6859 => x"38",
          6860 => x"2a",
          6861 => x"83",
          6862 => x"51",
          6863 => x"ff",
          6864 => x"b8",
          6865 => x"11",
          6866 => x"33",
          6867 => x"07",
          6868 => x"5a",
          6869 => x"ff",
          6870 => x"80",
          6871 => x"38",
          6872 => x"10",
          6873 => x"81",
          6874 => x"88",
          6875 => x"81",
          6876 => x"79",
          6877 => x"ff",
          6878 => x"7a",
          6879 => x"5c",
          6880 => x"72",
          6881 => x"38",
          6882 => x"85",
          6883 => x"55",
          6884 => x"33",
          6885 => x"71",
          6886 => x"57",
          6887 => x"38",
          6888 => x"ff",
          6889 => x"77",
          6890 => x"80",
          6891 => x"78",
          6892 => x"81",
          6893 => x"88",
          6894 => x"81",
          6895 => x"56",
          6896 => x"59",
          6897 => x"2e",
          6898 => x"59",
          6899 => x"73",
          6900 => x"38",
          6901 => x"80",
          6902 => x"38",
          6903 => x"82",
          6904 => x"16",
          6905 => x"78",
          6906 => x"80",
          6907 => x"88",
          6908 => x"56",
          6909 => x"74",
          6910 => x"15",
          6911 => x"d4",
          6912 => x"88",
          6913 => x"71",
          6914 => x"75",
          6915 => x"84",
          6916 => x"70",
          6917 => x"81",
          6918 => x"88",
          6919 => x"83",
          6920 => x"f8",
          6921 => x"7e",
          6922 => x"06",
          6923 => x"5c",
          6924 => x"59",
          6925 => x"82",
          6926 => x"81",
          6927 => x"72",
          6928 => x"84",
          6929 => x"18",
          6930 => x"34",
          6931 => x"34",
          6932 => x"08",
          6933 => x"11",
          6934 => x"33",
          6935 => x"71",
          6936 => x"74",
          6937 => x"5c",
          6938 => x"84",
          6939 => x"85",
          6940 => x"b8",
          6941 => x"16",
          6942 => x"86",
          6943 => x"12",
          6944 => x"2b",
          6945 => x"2a",
          6946 => x"59",
          6947 => x"34",
          6948 => x"34",
          6949 => x"08",
          6950 => x"11",
          6951 => x"33",
          6952 => x"71",
          6953 => x"74",
          6954 => x"5c",
          6955 => x"86",
          6956 => x"87",
          6957 => x"b8",
          6958 => x"16",
          6959 => x"84",
          6960 => x"12",
          6961 => x"2b",
          6962 => x"2a",
          6963 => x"59",
          6964 => x"34",
          6965 => x"34",
          6966 => x"08",
          6967 => x"51",
          6968 => x"e4",
          6969 => x"0d",
          6970 => x"33",
          6971 => x"71",
          6972 => x"83",
          6973 => x"05",
          6974 => x"85",
          6975 => x"88",
          6976 => x"88",
          6977 => x"59",
          6978 => x"74",
          6979 => x"76",
          6980 => x"84",
          6981 => x"70",
          6982 => x"33",
          6983 => x"71",
          6984 => x"83",
          6985 => x"05",
          6986 => x"87",
          6987 => x"88",
          6988 => x"88",
          6989 => x"5f",
          6990 => x"57",
          6991 => x"1a",
          6992 => x"1a",
          6993 => x"d4",
          6994 => x"33",
          6995 => x"71",
          6996 => x"81",
          6997 => x"70",
          6998 => x"57",
          6999 => x"77",
          7000 => x"18",
          7001 => x"d4",
          7002 => x"05",
          7003 => x"39",
          7004 => x"79",
          7005 => x"08",
          7006 => x"80",
          7007 => x"77",
          7008 => x"38",
          7009 => x"e4",
          7010 => x"0d",
          7011 => x"fb",
          7012 => x"b8",
          7013 => x"b8",
          7014 => x"3d",
          7015 => x"ff",
          7016 => x"b8",
          7017 => x"80",
          7018 => x"d0",
          7019 => x"80",
          7020 => x"84",
          7021 => x"fe",
          7022 => x"84",
          7023 => x"55",
          7024 => x"81",
          7025 => x"34",
          7026 => x"08",
          7027 => x"15",
          7028 => x"85",
          7029 => x"b8",
          7030 => x"76",
          7031 => x"81",
          7032 => x"34",
          7033 => x"08",
          7034 => x"22",
          7035 => x"80",
          7036 => x"83",
          7037 => x"70",
          7038 => x"51",
          7039 => x"88",
          7040 => x"89",
          7041 => x"b8",
          7042 => x"10",
          7043 => x"b8",
          7044 => x"f8",
          7045 => x"76",
          7046 => x"81",
          7047 => x"34",
          7048 => x"80",
          7049 => x"38",
          7050 => x"ed",
          7051 => x"67",
          7052 => x"70",
          7053 => x"08",
          7054 => x"76",
          7055 => x"aa",
          7056 => x"2e",
          7057 => x"7f",
          7058 => x"d7",
          7059 => x"84",
          7060 => x"38",
          7061 => x"83",
          7062 => x"70",
          7063 => x"06",
          7064 => x"83",
          7065 => x"7f",
          7066 => x"2a",
          7067 => x"ff",
          7068 => x"2b",
          7069 => x"33",
          7070 => x"71",
          7071 => x"70",
          7072 => x"83",
          7073 => x"70",
          7074 => x"fc",
          7075 => x"2b",
          7076 => x"33",
          7077 => x"71",
          7078 => x"70",
          7079 => x"90",
          7080 => x"45",
          7081 => x"54",
          7082 => x"48",
          7083 => x"5f",
          7084 => x"24",
          7085 => x"82",
          7086 => x"16",
          7087 => x"2b",
          7088 => x"10",
          7089 => x"33",
          7090 => x"71",
          7091 => x"90",
          7092 => x"5c",
          7093 => x"56",
          7094 => x"85",
          7095 => x"62",
          7096 => x"38",
          7097 => x"77",
          7098 => x"a2",
          7099 => x"2e",
          7100 => x"60",
          7101 => x"62",
          7102 => x"38",
          7103 => x"61",
          7104 => x"f7",
          7105 => x"70",
          7106 => x"33",
          7107 => x"71",
          7108 => x"7a",
          7109 => x"81",
          7110 => x"98",
          7111 => x"2b",
          7112 => x"59",
          7113 => x"5b",
          7114 => x"24",
          7115 => x"76",
          7116 => x"33",
          7117 => x"71",
          7118 => x"83",
          7119 => x"11",
          7120 => x"87",
          7121 => x"8b",
          7122 => x"2b",
          7123 => x"84",
          7124 => x"15",
          7125 => x"2b",
          7126 => x"2a",
          7127 => x"52",
          7128 => x"53",
          7129 => x"77",
          7130 => x"79",
          7131 => x"84",
          7132 => x"70",
          7133 => x"33",
          7134 => x"71",
          7135 => x"83",
          7136 => x"05",
          7137 => x"87",
          7138 => x"88",
          7139 => x"88",
          7140 => x"5e",
          7141 => x"41",
          7142 => x"16",
          7143 => x"16",
          7144 => x"d4",
          7145 => x"33",
          7146 => x"71",
          7147 => x"81",
          7148 => x"70",
          7149 => x"5c",
          7150 => x"79",
          7151 => x"1a",
          7152 => x"d4",
          7153 => x"82",
          7154 => x"12",
          7155 => x"2b",
          7156 => x"07",
          7157 => x"33",
          7158 => x"71",
          7159 => x"70",
          7160 => x"5c",
          7161 => x"5a",
          7162 => x"79",
          7163 => x"1a",
          7164 => x"d4",
          7165 => x"70",
          7166 => x"33",
          7167 => x"71",
          7168 => x"74",
          7169 => x"33",
          7170 => x"71",
          7171 => x"70",
          7172 => x"5c",
          7173 => x"5a",
          7174 => x"82",
          7175 => x"83",
          7176 => x"b8",
          7177 => x"1f",
          7178 => x"83",
          7179 => x"88",
          7180 => x"57",
          7181 => x"83",
          7182 => x"5a",
          7183 => x"84",
          7184 => x"c4",
          7185 => x"b8",
          7186 => x"84",
          7187 => x"05",
          7188 => x"ff",
          7189 => x"44",
          7190 => x"26",
          7191 => x"7e",
          7192 => x"b8",
          7193 => x"3d",
          7194 => x"ff",
          7195 => x"b8",
          7196 => x"80",
          7197 => x"d0",
          7198 => x"80",
          7199 => x"84",
          7200 => x"fe",
          7201 => x"84",
          7202 => x"5e",
          7203 => x"81",
          7204 => x"34",
          7205 => x"08",
          7206 => x"1e",
          7207 => x"85",
          7208 => x"b8",
          7209 => x"60",
          7210 => x"81",
          7211 => x"34",
          7212 => x"08",
          7213 => x"22",
          7214 => x"80",
          7215 => x"83",
          7216 => x"70",
          7217 => x"5a",
          7218 => x"88",
          7219 => x"89",
          7220 => x"b8",
          7221 => x"10",
          7222 => x"b8",
          7223 => x"f8",
          7224 => x"60",
          7225 => x"81",
          7226 => x"34",
          7227 => x"08",
          7228 => x"d3",
          7229 => x"2e",
          7230 => x"7e",
          7231 => x"2e",
          7232 => x"7f",
          7233 => x"3f",
          7234 => x"08",
          7235 => x"0c",
          7236 => x"04",
          7237 => x"b8",
          7238 => x"83",
          7239 => x"5e",
          7240 => x"70",
          7241 => x"33",
          7242 => x"07",
          7243 => x"06",
          7244 => x"48",
          7245 => x"40",
          7246 => x"60",
          7247 => x"61",
          7248 => x"08",
          7249 => x"2a",
          7250 => x"82",
          7251 => x"83",
          7252 => x"b8",
          7253 => x"1f",
          7254 => x"12",
          7255 => x"2b",
          7256 => x"2b",
          7257 => x"06",
          7258 => x"83",
          7259 => x"70",
          7260 => x"5c",
          7261 => x"5b",
          7262 => x"82",
          7263 => x"81",
          7264 => x"60",
          7265 => x"34",
          7266 => x"08",
          7267 => x"7b",
          7268 => x"1c",
          7269 => x"b8",
          7270 => x"84",
          7271 => x"88",
          7272 => x"fd",
          7273 => x"75",
          7274 => x"ff",
          7275 => x"54",
          7276 => x"77",
          7277 => x"06",
          7278 => x"83",
          7279 => x"82",
          7280 => x"18",
          7281 => x"2b",
          7282 => x"10",
          7283 => x"33",
          7284 => x"71",
          7285 => x"90",
          7286 => x"5e",
          7287 => x"58",
          7288 => x"80",
          7289 => x"38",
          7290 => x"61",
          7291 => x"83",
          7292 => x"24",
          7293 => x"77",
          7294 => x"06",
          7295 => x"27",
          7296 => x"fe",
          7297 => x"ff",
          7298 => x"b8",
          7299 => x"80",
          7300 => x"d0",
          7301 => x"80",
          7302 => x"84",
          7303 => x"fe",
          7304 => x"84",
          7305 => x"5a",
          7306 => x"81",
          7307 => x"34",
          7308 => x"08",
          7309 => x"1a",
          7310 => x"85",
          7311 => x"b8",
          7312 => x"7e",
          7313 => x"81",
          7314 => x"34",
          7315 => x"08",
          7316 => x"22",
          7317 => x"80",
          7318 => x"83",
          7319 => x"70",
          7320 => x"56",
          7321 => x"64",
          7322 => x"73",
          7323 => x"34",
          7324 => x"22",
          7325 => x"10",
          7326 => x"08",
          7327 => x"42",
          7328 => x"82",
          7329 => x"61",
          7330 => x"fc",
          7331 => x"7a",
          7332 => x"38",
          7333 => x"ff",
          7334 => x"7b",
          7335 => x"38",
          7336 => x"76",
          7337 => x"bd",
          7338 => x"ea",
          7339 => x"54",
          7340 => x"e4",
          7341 => x"0d",
          7342 => x"82",
          7343 => x"12",
          7344 => x"2b",
          7345 => x"07",
          7346 => x"11",
          7347 => x"33",
          7348 => x"71",
          7349 => x"7e",
          7350 => x"33",
          7351 => x"71",
          7352 => x"70",
          7353 => x"44",
          7354 => x"46",
          7355 => x"45",
          7356 => x"84",
          7357 => x"64",
          7358 => x"84",
          7359 => x"70",
          7360 => x"33",
          7361 => x"71",
          7362 => x"83",
          7363 => x"05",
          7364 => x"87",
          7365 => x"88",
          7366 => x"88",
          7367 => x"42",
          7368 => x"5d",
          7369 => x"86",
          7370 => x"64",
          7371 => x"84",
          7372 => x"16",
          7373 => x"12",
          7374 => x"2b",
          7375 => x"ff",
          7376 => x"2a",
          7377 => x"5d",
          7378 => x"79",
          7379 => x"84",
          7380 => x"70",
          7381 => x"33",
          7382 => x"71",
          7383 => x"83",
          7384 => x"05",
          7385 => x"15",
          7386 => x"2b",
          7387 => x"2a",
          7388 => x"40",
          7389 => x"54",
          7390 => x"75",
          7391 => x"84",
          7392 => x"70",
          7393 => x"81",
          7394 => x"8b",
          7395 => x"2b",
          7396 => x"82",
          7397 => x"15",
          7398 => x"2b",
          7399 => x"2a",
          7400 => x"5b",
          7401 => x"55",
          7402 => x"34",
          7403 => x"34",
          7404 => x"08",
          7405 => x"11",
          7406 => x"33",
          7407 => x"07",
          7408 => x"56",
          7409 => x"42",
          7410 => x"7e",
          7411 => x"51",
          7412 => x"3f",
          7413 => x"08",
          7414 => x"78",
          7415 => x"06",
          7416 => x"99",
          7417 => x"f4",
          7418 => x"d4",
          7419 => x"0b",
          7420 => x"23",
          7421 => x"53",
          7422 => x"ff",
          7423 => x"c0",
          7424 => x"b8",
          7425 => x"7f",
          7426 => x"0b",
          7427 => x"84",
          7428 => x"55",
          7429 => x"34",
          7430 => x"16",
          7431 => x"d4",
          7432 => x"86",
          7433 => x"0b",
          7434 => x"84",
          7435 => x"84",
          7436 => x"ff",
          7437 => x"80",
          7438 => x"ff",
          7439 => x"88",
          7440 => x"44",
          7441 => x"1f",
          7442 => x"1f",
          7443 => x"d0",
          7444 => x"10",
          7445 => x"d4",
          7446 => x"05",
          7447 => x"82",
          7448 => x"0b",
          7449 => x"7e",
          7450 => x"3f",
          7451 => x"c0",
          7452 => x"33",
          7453 => x"71",
          7454 => x"83",
          7455 => x"05",
          7456 => x"85",
          7457 => x"88",
          7458 => x"88",
          7459 => x"5e",
          7460 => x"76",
          7461 => x"34",
          7462 => x"05",
          7463 => x"d4",
          7464 => x"84",
          7465 => x"12",
          7466 => x"2b",
          7467 => x"07",
          7468 => x"14",
          7469 => x"33",
          7470 => x"07",
          7471 => x"41",
          7472 => x"59",
          7473 => x"79",
          7474 => x"34",
          7475 => x"05",
          7476 => x"d4",
          7477 => x"33",
          7478 => x"71",
          7479 => x"81",
          7480 => x"70",
          7481 => x"42",
          7482 => x"78",
          7483 => x"19",
          7484 => x"d4",
          7485 => x"70",
          7486 => x"33",
          7487 => x"71",
          7488 => x"74",
          7489 => x"81",
          7490 => x"88",
          7491 => x"83",
          7492 => x"f8",
          7493 => x"63",
          7494 => x"5d",
          7495 => x"40",
          7496 => x"7f",
          7497 => x"7b",
          7498 => x"84",
          7499 => x"70",
          7500 => x"81",
          7501 => x"8b",
          7502 => x"2b",
          7503 => x"70",
          7504 => x"33",
          7505 => x"07",
          7506 => x"06",
          7507 => x"48",
          7508 => x"46",
          7509 => x"60",
          7510 => x"60",
          7511 => x"61",
          7512 => x"06",
          7513 => x"39",
          7514 => x"87",
          7515 => x"8b",
          7516 => x"2b",
          7517 => x"84",
          7518 => x"19",
          7519 => x"2b",
          7520 => x"2a",
          7521 => x"52",
          7522 => x"84",
          7523 => x"85",
          7524 => x"b8",
          7525 => x"19",
          7526 => x"85",
          7527 => x"8b",
          7528 => x"2b",
          7529 => x"86",
          7530 => x"15",
          7531 => x"2b",
          7532 => x"2a",
          7533 => x"52",
          7534 => x"56",
          7535 => x"05",
          7536 => x"87",
          7537 => x"b8",
          7538 => x"70",
          7539 => x"33",
          7540 => x"07",
          7541 => x"06",
          7542 => x"5b",
          7543 => x"77",
          7544 => x"81",
          7545 => x"b8",
          7546 => x"1f",
          7547 => x"12",
          7548 => x"2b",
          7549 => x"07",
          7550 => x"33",
          7551 => x"71",
          7552 => x"70",
          7553 => x"ff",
          7554 => x"05",
          7555 => x"56",
          7556 => x"58",
          7557 => x"55",
          7558 => x"34",
          7559 => x"34",
          7560 => x"08",
          7561 => x"33",
          7562 => x"71",
          7563 => x"83",
          7564 => x"05",
          7565 => x"12",
          7566 => x"2b",
          7567 => x"ff",
          7568 => x"2a",
          7569 => x"58",
          7570 => x"55",
          7571 => x"76",
          7572 => x"84",
          7573 => x"70",
          7574 => x"33",
          7575 => x"71",
          7576 => x"83",
          7577 => x"11",
          7578 => x"87",
          7579 => x"8b",
          7580 => x"2b",
          7581 => x"84",
          7582 => x"15",
          7583 => x"2b",
          7584 => x"2a",
          7585 => x"52",
          7586 => x"53",
          7587 => x"57",
          7588 => x"34",
          7589 => x"34",
          7590 => x"08",
          7591 => x"11",
          7592 => x"33",
          7593 => x"71",
          7594 => x"74",
          7595 => x"33",
          7596 => x"71",
          7597 => x"70",
          7598 => x"42",
          7599 => x"57",
          7600 => x"86",
          7601 => x"87",
          7602 => x"b8",
          7603 => x"70",
          7604 => x"33",
          7605 => x"07",
          7606 => x"06",
          7607 => x"5a",
          7608 => x"76",
          7609 => x"81",
          7610 => x"b8",
          7611 => x"1f",
          7612 => x"83",
          7613 => x"8b",
          7614 => x"2b",
          7615 => x"73",
          7616 => x"33",
          7617 => x"07",
          7618 => x"41",
          7619 => x"5f",
          7620 => x"79",
          7621 => x"81",
          7622 => x"b8",
          7623 => x"1f",
          7624 => x"12",
          7625 => x"2b",
          7626 => x"07",
          7627 => x"14",
          7628 => x"33",
          7629 => x"07",
          7630 => x"41",
          7631 => x"5f",
          7632 => x"79",
          7633 => x"75",
          7634 => x"84",
          7635 => x"70",
          7636 => x"33",
          7637 => x"71",
          7638 => x"66",
          7639 => x"70",
          7640 => x"52",
          7641 => x"05",
          7642 => x"fe",
          7643 => x"84",
          7644 => x"1e",
          7645 => x"65",
          7646 => x"83",
          7647 => x"5d",
          7648 => x"d5",
          7649 => x"33",
          7650 => x"71",
          7651 => x"83",
          7652 => x"05",
          7653 => x"85",
          7654 => x"88",
          7655 => x"88",
          7656 => x"5d",
          7657 => x"7a",
          7658 => x"34",
          7659 => x"05",
          7660 => x"d4",
          7661 => x"84",
          7662 => x"12",
          7663 => x"2b",
          7664 => x"07",
          7665 => x"14",
          7666 => x"33",
          7667 => x"07",
          7668 => x"5b",
          7669 => x"5c",
          7670 => x"73",
          7671 => x"34",
          7672 => x"05",
          7673 => x"d4",
          7674 => x"33",
          7675 => x"71",
          7676 => x"81",
          7677 => x"70",
          7678 => x"5f",
          7679 => x"75",
          7680 => x"16",
          7681 => x"d4",
          7682 => x"70",
          7683 => x"33",
          7684 => x"71",
          7685 => x"74",
          7686 => x"81",
          7687 => x"88",
          7688 => x"83",
          7689 => x"f8",
          7690 => x"63",
          7691 => x"44",
          7692 => x"5e",
          7693 => x"74",
          7694 => x"7b",
          7695 => x"84",
          7696 => x"70",
          7697 => x"81",
          7698 => x"8b",
          7699 => x"2b",
          7700 => x"70",
          7701 => x"33",
          7702 => x"07",
          7703 => x"06",
          7704 => x"47",
          7705 => x"46",
          7706 => x"7f",
          7707 => x"81",
          7708 => x"83",
          7709 => x"5b",
          7710 => x"7e",
          7711 => x"e5",
          7712 => x"b8",
          7713 => x"84",
          7714 => x"80",
          7715 => x"62",
          7716 => x"84",
          7717 => x"51",
          7718 => x"3f",
          7719 => x"88",
          7720 => x"61",
          7721 => x"b7",
          7722 => x"39",
          7723 => x"7a",
          7724 => x"b8",
          7725 => x"58",
          7726 => x"b7",
          7727 => x"77",
          7728 => x"84",
          7729 => x"89",
          7730 => x"77",
          7731 => x"3f",
          7732 => x"08",
          7733 => x"e4",
          7734 => x"e6",
          7735 => x"80",
          7736 => x"e4",
          7737 => x"b7",
          7738 => x"84",
          7739 => x"89",
          7740 => x"84",
          7741 => x"84",
          7742 => x"a0",
          7743 => x"b8",
          7744 => x"80",
          7745 => x"52",
          7746 => x"51",
          7747 => x"3f",
          7748 => x"08",
          7749 => x"34",
          7750 => x"16",
          7751 => x"d4",
          7752 => x"84",
          7753 => x"0b",
          7754 => x"84",
          7755 => x"56",
          7756 => x"34",
          7757 => x"17",
          7758 => x"d4",
          7759 => x"d0",
          7760 => x"fe",
          7761 => x"70",
          7762 => x"06",
          7763 => x"58",
          7764 => x"74",
          7765 => x"73",
          7766 => x"84",
          7767 => x"70",
          7768 => x"84",
          7769 => x"05",
          7770 => x"55",
          7771 => x"34",
          7772 => x"15",
          7773 => x"77",
          7774 => x"c6",
          7775 => x"39",
          7776 => x"02",
          7777 => x"51",
          7778 => x"72",
          7779 => x"84",
          7780 => x"33",
          7781 => x"b8",
          7782 => x"3d",
          7783 => x"3d",
          7784 => x"05",
          7785 => x"53",
          7786 => x"9d",
          7787 => x"d4",
          7788 => x"b8",
          7789 => x"ff",
          7790 => x"87",
          7791 => x"b8",
          7792 => x"84",
          7793 => x"33",
          7794 => x"b8",
          7795 => x"3d",
          7796 => x"3d",
          7797 => x"60",
          7798 => x"af",
          7799 => x"5c",
          7800 => x"54",
          7801 => x"87",
          7802 => x"e0",
          7803 => x"73",
          7804 => x"83",
          7805 => x"38",
          7806 => x"0b",
          7807 => x"8c",
          7808 => x"75",
          7809 => x"d5",
          7810 => x"b8",
          7811 => x"ff",
          7812 => x"80",
          7813 => x"87",
          7814 => x"08",
          7815 => x"38",
          7816 => x"d6",
          7817 => x"80",
          7818 => x"73",
          7819 => x"38",
          7820 => x"55",
          7821 => x"e4",
          7822 => x"0d",
          7823 => x"16",
          7824 => x"81",
          7825 => x"55",
          7826 => x"26",
          7827 => x"d5",
          7828 => x"0d",
          7829 => x"02",
          7830 => x"05",
          7831 => x"57",
          7832 => x"76",
          7833 => x"38",
          7834 => x"17",
          7835 => x"81",
          7836 => x"55",
          7837 => x"73",
          7838 => x"87",
          7839 => x"0c",
          7840 => x"52",
          7841 => x"8e",
          7842 => x"e4",
          7843 => x"06",
          7844 => x"2e",
          7845 => x"c0",
          7846 => x"54",
          7847 => x"79",
          7848 => x"38",
          7849 => x"80",
          7850 => x"80",
          7851 => x"81",
          7852 => x"74",
          7853 => x"0c",
          7854 => x"04",
          7855 => x"81",
          7856 => x"ff",
          7857 => x"56",
          7858 => x"ff",
          7859 => x"39",
          7860 => x"78",
          7861 => x"9b",
          7862 => x"88",
          7863 => x"33",
          7864 => x"81",
          7865 => x"26",
          7866 => x"b8",
          7867 => x"53",
          7868 => x"54",
          7869 => x"9b",
          7870 => x"87",
          7871 => x"0c",
          7872 => x"73",
          7873 => x"72",
          7874 => x"38",
          7875 => x"9a",
          7876 => x"72",
          7877 => x"0c",
          7878 => x"04",
          7879 => x"75",
          7880 => x"b8",
          7881 => x"3d",
          7882 => x"80",
          7883 => x"0b",
          7884 => x"0c",
          7885 => x"04",
          7886 => x"87",
          7887 => x"11",
          7888 => x"cd",
          7889 => x"70",
          7890 => x"06",
          7891 => x"80",
          7892 => x"87",
          7893 => x"08",
          7894 => x"38",
          7895 => x"8c",
          7896 => x"ca",
          7897 => x"0c",
          7898 => x"8c",
          7899 => x"08",
          7900 => x"73",
          7901 => x"9b",
          7902 => x"82",
          7903 => x"ee",
          7904 => x"39",
          7905 => x"7c",
          7906 => x"83",
          7907 => x"5b",
          7908 => x"77",
          7909 => x"06",
          7910 => x"33",
          7911 => x"2e",
          7912 => x"80",
          7913 => x"81",
          7914 => x"fe",
          7915 => x"b8",
          7916 => x"2e",
          7917 => x"59",
          7918 => x"e4",
          7919 => x"0d",
          7920 => x"b4",
          7921 => x"b8",
          7922 => x"81",
          7923 => x"5a",
          7924 => x"81",
          7925 => x"e4",
          7926 => x"09",
          7927 => x"38",
          7928 => x"08",
          7929 => x"b4",
          7930 => x"a8",
          7931 => x"a0",
          7932 => x"b8",
          7933 => x"58",
          7934 => x"76",
          7935 => x"38",
          7936 => x"55",
          7937 => x"09",
          7938 => x"8e",
          7939 => x"75",
          7940 => x"52",
          7941 => x"51",
          7942 => x"76",
          7943 => x"59",
          7944 => x"09",
          7945 => x"fb",
          7946 => x"33",
          7947 => x"2e",
          7948 => x"fe",
          7949 => x"18",
          7950 => x"7a",
          7951 => x"75",
          7952 => x"57",
          7953 => x"57",
          7954 => x"80",
          7955 => x"b6",
          7956 => x"aa",
          7957 => x"19",
          7958 => x"7a",
          7959 => x"0b",
          7960 => x"80",
          7961 => x"19",
          7962 => x"0b",
          7963 => x"80",
          7964 => x"9c",
          7965 => x"f2",
          7966 => x"19",
          7967 => x"0b",
          7968 => x"34",
          7969 => x"84",
          7970 => x"94",
          7971 => x"74",
          7972 => x"34",
          7973 => x"5b",
          7974 => x"19",
          7975 => x"2a",
          7976 => x"a2",
          7977 => x"98",
          7978 => x"84",
          7979 => x"90",
          7980 => x"7a",
          7981 => x"34",
          7982 => x"55",
          7983 => x"19",
          7984 => x"2a",
          7985 => x"a6",
          7986 => x"98",
          7987 => x"84",
          7988 => x"a4",
          7989 => x"05",
          7990 => x"0c",
          7991 => x"7a",
          7992 => x"81",
          7993 => x"fa",
          7994 => x"84",
          7995 => x"53",
          7996 => x"18",
          7997 => x"d8",
          7998 => x"e4",
          7999 => x"fd",
          8000 => x"b2",
          8001 => x"0d",
          8002 => x"08",
          8003 => x"81",
          8004 => x"38",
          8005 => x"76",
          8006 => x"81",
          8007 => x"b8",
          8008 => x"3d",
          8009 => x"77",
          8010 => x"74",
          8011 => x"cc",
          8012 => x"24",
          8013 => x"74",
          8014 => x"81",
          8015 => x"75",
          8016 => x"70",
          8017 => x"19",
          8018 => x"5a",
          8019 => x"17",
          8020 => x"b0",
          8021 => x"33",
          8022 => x"2e",
          8023 => x"83",
          8024 => x"54",
          8025 => x"17",
          8026 => x"33",
          8027 => x"3f",
          8028 => x"08",
          8029 => x"38",
          8030 => x"5b",
          8031 => x"0c",
          8032 => x"38",
          8033 => x"06",
          8034 => x"33",
          8035 => x"89",
          8036 => x"08",
          8037 => x"5d",
          8038 => x"08",
          8039 => x"38",
          8040 => x"18",
          8041 => x"56",
          8042 => x"2e",
          8043 => x"84",
          8044 => x"54",
          8045 => x"17",
          8046 => x"33",
          8047 => x"3f",
          8048 => x"08",
          8049 => x"38",
          8050 => x"5a",
          8051 => x"0c",
          8052 => x"38",
          8053 => x"06",
          8054 => x"33",
          8055 => x"7e",
          8056 => x"06",
          8057 => x"53",
          8058 => x"5d",
          8059 => x"38",
          8060 => x"06",
          8061 => x"0c",
          8062 => x"04",
          8063 => x"a8",
          8064 => x"59",
          8065 => x"79",
          8066 => x"80",
          8067 => x"33",
          8068 => x"5b",
          8069 => x"09",
          8070 => x"c2",
          8071 => x"78",
          8072 => x"52",
          8073 => x"51",
          8074 => x"84",
          8075 => x"80",
          8076 => x"ff",
          8077 => x"78",
          8078 => x"79",
          8079 => x"75",
          8080 => x"06",
          8081 => x"05",
          8082 => x"71",
          8083 => x"2b",
          8084 => x"e4",
          8085 => x"8f",
          8086 => x"74",
          8087 => x"81",
          8088 => x"38",
          8089 => x"a8",
          8090 => x"59",
          8091 => x"79",
          8092 => x"80",
          8093 => x"33",
          8094 => x"5b",
          8095 => x"09",
          8096 => x"81",
          8097 => x"78",
          8098 => x"52",
          8099 => x"51",
          8100 => x"84",
          8101 => x"80",
          8102 => x"ff",
          8103 => x"78",
          8104 => x"79",
          8105 => x"75",
          8106 => x"fc",
          8107 => x"b8",
          8108 => x"33",
          8109 => x"71",
          8110 => x"88",
          8111 => x"14",
          8112 => x"07",
          8113 => x"33",
          8114 => x"ff",
          8115 => x"07",
          8116 => x"0c",
          8117 => x"59",
          8118 => x"3d",
          8119 => x"54",
          8120 => x"53",
          8121 => x"53",
          8122 => x"52",
          8123 => x"3f",
          8124 => x"b8",
          8125 => x"2e",
          8126 => x"fe",
          8127 => x"b8",
          8128 => x"18",
          8129 => x"08",
          8130 => x"31",
          8131 => x"08",
          8132 => x"a0",
          8133 => x"fe",
          8134 => x"17",
          8135 => x"82",
          8136 => x"06",
          8137 => x"81",
          8138 => x"08",
          8139 => x"05",
          8140 => x"81",
          8141 => x"f6",
          8142 => x"5a",
          8143 => x"81",
          8144 => x"08",
          8145 => x"70",
          8146 => x"33",
          8147 => x"81",
          8148 => x"e4",
          8149 => x"09",
          8150 => x"81",
          8151 => x"e4",
          8152 => x"34",
          8153 => x"a8",
          8154 => x"5d",
          8155 => x"08",
          8156 => x"82",
          8157 => x"7d",
          8158 => x"cb",
          8159 => x"e4",
          8160 => x"de",
          8161 => x"b4",
          8162 => x"b8",
          8163 => x"81",
          8164 => x"5c",
          8165 => x"81",
          8166 => x"e4",
          8167 => x"09",
          8168 => x"ff",
          8169 => x"e4",
          8170 => x"34",
          8171 => x"a8",
          8172 => x"84",
          8173 => x"5b",
          8174 => x"18",
          8175 => x"c5",
          8176 => x"33",
          8177 => x"2e",
          8178 => x"fd",
          8179 => x"54",
          8180 => x"a0",
          8181 => x"53",
          8182 => x"17",
          8183 => x"f1",
          8184 => x"fd",
          8185 => x"54",
          8186 => x"53",
          8187 => x"53",
          8188 => x"52",
          8189 => x"3f",
          8190 => x"b8",
          8191 => x"2e",
          8192 => x"fb",
          8193 => x"b8",
          8194 => x"18",
          8195 => x"08",
          8196 => x"31",
          8197 => x"08",
          8198 => x"a0",
          8199 => x"fb",
          8200 => x"17",
          8201 => x"82",
          8202 => x"06",
          8203 => x"81",
          8204 => x"08",
          8205 => x"05",
          8206 => x"81",
          8207 => x"f4",
          8208 => x"5a",
          8209 => x"81",
          8210 => x"08",
          8211 => x"05",
          8212 => x"81",
          8213 => x"f3",
          8214 => x"86",
          8215 => x"7a",
          8216 => x"fa",
          8217 => x"3d",
          8218 => x"64",
          8219 => x"82",
          8220 => x"27",
          8221 => x"9c",
          8222 => x"95",
          8223 => x"55",
          8224 => x"96",
          8225 => x"24",
          8226 => x"74",
          8227 => x"8a",
          8228 => x"b8",
          8229 => x"3d",
          8230 => x"88",
          8231 => x"08",
          8232 => x"0b",
          8233 => x"58",
          8234 => x"2e",
          8235 => x"83",
          8236 => x"5b",
          8237 => x"2e",
          8238 => x"83",
          8239 => x"54",
          8240 => x"19",
          8241 => x"33",
          8242 => x"3f",
          8243 => x"08",
          8244 => x"38",
          8245 => x"5a",
          8246 => x"0c",
          8247 => x"ff",
          8248 => x"10",
          8249 => x"79",
          8250 => x"ff",
          8251 => x"5e",
          8252 => x"34",
          8253 => x"5a",
          8254 => x"34",
          8255 => x"1a",
          8256 => x"b8",
          8257 => x"3d",
          8258 => x"83",
          8259 => x"06",
          8260 => x"75",
          8261 => x"1a",
          8262 => x"80",
          8263 => x"08",
          8264 => x"78",
          8265 => x"38",
          8266 => x"7c",
          8267 => x"7c",
          8268 => x"06",
          8269 => x"81",
          8270 => x"b8",
          8271 => x"19",
          8272 => x"8e",
          8273 => x"e4",
          8274 => x"85",
          8275 => x"81",
          8276 => x"1a",
          8277 => x"79",
          8278 => x"75",
          8279 => x"fc",
          8280 => x"b8",
          8281 => x"33",
          8282 => x"8f",
          8283 => x"f0",
          8284 => x"41",
          8285 => x"7d",
          8286 => x"88",
          8287 => x"b9",
          8288 => x"90",
          8289 => x"ba",
          8290 => x"98",
          8291 => x"bb",
          8292 => x"0b",
          8293 => x"fe",
          8294 => x"81",
          8295 => x"89",
          8296 => x"08",
          8297 => x"08",
          8298 => x"76",
          8299 => x"38",
          8300 => x"1a",
          8301 => x"56",
          8302 => x"2e",
          8303 => x"82",
          8304 => x"54",
          8305 => x"19",
          8306 => x"33",
          8307 => x"3f",
          8308 => x"08",
          8309 => x"38",
          8310 => x"5c",
          8311 => x"0c",
          8312 => x"fd",
          8313 => x"83",
          8314 => x"b8",
          8315 => x"77",
          8316 => x"5f",
          8317 => x"7c",
          8318 => x"38",
          8319 => x"9f",
          8320 => x"33",
          8321 => x"07",
          8322 => x"77",
          8323 => x"83",
          8324 => x"89",
          8325 => x"08",
          8326 => x"0b",
          8327 => x"56",
          8328 => x"2e",
          8329 => x"81",
          8330 => x"b8",
          8331 => x"81",
          8332 => x"57",
          8333 => x"81",
          8334 => x"e4",
          8335 => x"09",
          8336 => x"c7",
          8337 => x"e4",
          8338 => x"34",
          8339 => x"70",
          8340 => x"31",
          8341 => x"84",
          8342 => x"5b",
          8343 => x"74",
          8344 => x"38",
          8345 => x"55",
          8346 => x"82",
          8347 => x"54",
          8348 => x"52",
          8349 => x"51",
          8350 => x"84",
          8351 => x"80",
          8352 => x"ff",
          8353 => x"75",
          8354 => x"77",
          8355 => x"7d",
          8356 => x"19",
          8357 => x"84",
          8358 => x"7c",
          8359 => x"88",
          8360 => x"81",
          8361 => x"8f",
          8362 => x"5c",
          8363 => x"81",
          8364 => x"34",
          8365 => x"81",
          8366 => x"b8",
          8367 => x"81",
          8368 => x"5d",
          8369 => x"81",
          8370 => x"e4",
          8371 => x"09",
          8372 => x"88",
          8373 => x"e4",
          8374 => x"34",
          8375 => x"70",
          8376 => x"31",
          8377 => x"84",
          8378 => x"5d",
          8379 => x"7e",
          8380 => x"ca",
          8381 => x"33",
          8382 => x"2e",
          8383 => x"fb",
          8384 => x"54",
          8385 => x"7c",
          8386 => x"33",
          8387 => x"3f",
          8388 => x"aa",
          8389 => x"76",
          8390 => x"70",
          8391 => x"33",
          8392 => x"ad",
          8393 => x"84",
          8394 => x"7d",
          8395 => x"06",
          8396 => x"84",
          8397 => x"83",
          8398 => x"19",
          8399 => x"1b",
          8400 => x"1b",
          8401 => x"e4",
          8402 => x"56",
          8403 => x"27",
          8404 => x"82",
          8405 => x"74",
          8406 => x"81",
          8407 => x"38",
          8408 => x"1f",
          8409 => x"81",
          8410 => x"ed",
          8411 => x"5c",
          8412 => x"81",
          8413 => x"b8",
          8414 => x"81",
          8415 => x"57",
          8416 => x"81",
          8417 => x"e4",
          8418 => x"09",
          8419 => x"c5",
          8420 => x"e4",
          8421 => x"34",
          8422 => x"70",
          8423 => x"31",
          8424 => x"84",
          8425 => x"5d",
          8426 => x"7e",
          8427 => x"87",
          8428 => x"33",
          8429 => x"2e",
          8430 => x"fa",
          8431 => x"54",
          8432 => x"76",
          8433 => x"33",
          8434 => x"3f",
          8435 => x"e7",
          8436 => x"79",
          8437 => x"52",
          8438 => x"51",
          8439 => x"7e",
          8440 => x"39",
          8441 => x"83",
          8442 => x"05",
          8443 => x"ff",
          8444 => x"58",
          8445 => x"34",
          8446 => x"5a",
          8447 => x"34",
          8448 => x"7e",
          8449 => x"39",
          8450 => x"2b",
          8451 => x"7a",
          8452 => x"83",
          8453 => x"98",
          8454 => x"06",
          8455 => x"06",
          8456 => x"5f",
          8457 => x"7d",
          8458 => x"2a",
          8459 => x"1d",
          8460 => x"2a",
          8461 => x"1d",
          8462 => x"2a",
          8463 => x"1d",
          8464 => x"39",
          8465 => x"7c",
          8466 => x"5b",
          8467 => x"81",
          8468 => x"19",
          8469 => x"80",
          8470 => x"38",
          8471 => x"08",
          8472 => x"38",
          8473 => x"70",
          8474 => x"80",
          8475 => x"38",
          8476 => x"81",
          8477 => x"56",
          8478 => x"9c",
          8479 => x"26",
          8480 => x"56",
          8481 => x"82",
          8482 => x"52",
          8483 => x"f5",
          8484 => x"e4",
          8485 => x"81",
          8486 => x"58",
          8487 => x"08",
          8488 => x"38",
          8489 => x"08",
          8490 => x"70",
          8491 => x"25",
          8492 => x"51",
          8493 => x"73",
          8494 => x"75",
          8495 => x"81",
          8496 => x"38",
          8497 => x"84",
          8498 => x"8c",
          8499 => x"81",
          8500 => x"39",
          8501 => x"08",
          8502 => x"7a",
          8503 => x"f0",
          8504 => x"55",
          8505 => x"e4",
          8506 => x"38",
          8507 => x"08",
          8508 => x"e4",
          8509 => x"ce",
          8510 => x"08",
          8511 => x"08",
          8512 => x"7a",
          8513 => x"39",
          8514 => x"9c",
          8515 => x"26",
          8516 => x"56",
          8517 => x"51",
          8518 => x"80",
          8519 => x"e4",
          8520 => x"81",
          8521 => x"b8",
          8522 => x"70",
          8523 => x"07",
          8524 => x"7b",
          8525 => x"e4",
          8526 => x"51",
          8527 => x"ff",
          8528 => x"b8",
          8529 => x"2e",
          8530 => x"19",
          8531 => x"74",
          8532 => x"38",
          8533 => x"08",
          8534 => x"38",
          8535 => x"57",
          8536 => x"75",
          8537 => x"8e",
          8538 => x"75",
          8539 => x"f5",
          8540 => x"b8",
          8541 => x"b8",
          8542 => x"70",
          8543 => x"08",
          8544 => x"56",
          8545 => x"80",
          8546 => x"80",
          8547 => x"90",
          8548 => x"19",
          8549 => x"94",
          8550 => x"58",
          8551 => x"86",
          8552 => x"94",
          8553 => x"19",
          8554 => x"5a",
          8555 => x"34",
          8556 => x"84",
          8557 => x"8c",
          8558 => x"80",
          8559 => x"e4",
          8560 => x"0d",
          8561 => x"e4",
          8562 => x"da",
          8563 => x"2e",
          8564 => x"75",
          8565 => x"78",
          8566 => x"3f",
          8567 => x"08",
          8568 => x"39",
          8569 => x"08",
          8570 => x"0c",
          8571 => x"04",
          8572 => x"81",
          8573 => x"38",
          8574 => x"b6",
          8575 => x"0d",
          8576 => x"08",
          8577 => x"73",
          8578 => x"26",
          8579 => x"73",
          8580 => x"72",
          8581 => x"73",
          8582 => x"88",
          8583 => x"74",
          8584 => x"76",
          8585 => x"82",
          8586 => x"38",
          8587 => x"53",
          8588 => x"18",
          8589 => x"72",
          8590 => x"38",
          8591 => x"98",
          8592 => x"94",
          8593 => x"18",
          8594 => x"56",
          8595 => x"94",
          8596 => x"2a",
          8597 => x"0c",
          8598 => x"06",
          8599 => x"9c",
          8600 => x"56",
          8601 => x"e4",
          8602 => x"0d",
          8603 => x"84",
          8604 => x"8a",
          8605 => x"ac",
          8606 => x"74",
          8607 => x"ac",
          8608 => x"22",
          8609 => x"57",
          8610 => x"27",
          8611 => x"17",
          8612 => x"15",
          8613 => x"56",
          8614 => x"73",
          8615 => x"8a",
          8616 => x"71",
          8617 => x"08",
          8618 => x"78",
          8619 => x"ff",
          8620 => x"52",
          8621 => x"cd",
          8622 => x"e4",
          8623 => x"b8",
          8624 => x"2e",
          8625 => x"0b",
          8626 => x"08",
          8627 => x"38",
          8628 => x"53",
          8629 => x"08",
          8630 => x"91",
          8631 => x"31",
          8632 => x"27",
          8633 => x"aa",
          8634 => x"84",
          8635 => x"8a",
          8636 => x"f3",
          8637 => x"70",
          8638 => x"08",
          8639 => x"5a",
          8640 => x"0a",
          8641 => x"38",
          8642 => x"18",
          8643 => x"08",
          8644 => x"74",
          8645 => x"38",
          8646 => x"06",
          8647 => x"38",
          8648 => x"18",
          8649 => x"75",
          8650 => x"85",
          8651 => x"22",
          8652 => x"76",
          8653 => x"38",
          8654 => x"0c",
          8655 => x"0c",
          8656 => x"05",
          8657 => x"80",
          8658 => x"b8",
          8659 => x"3d",
          8660 => x"98",
          8661 => x"19",
          8662 => x"7a",
          8663 => x"5c",
          8664 => x"75",
          8665 => x"eb",
          8666 => x"b8",
          8667 => x"82",
          8668 => x"84",
          8669 => x"27",
          8670 => x"56",
          8671 => x"08",
          8672 => x"38",
          8673 => x"84",
          8674 => x"26",
          8675 => x"60",
          8676 => x"98",
          8677 => x"08",
          8678 => x"f9",
          8679 => x"b8",
          8680 => x"87",
          8681 => x"e4",
          8682 => x"ff",
          8683 => x"56",
          8684 => x"08",
          8685 => x"91",
          8686 => x"84",
          8687 => x"ff",
          8688 => x"38",
          8689 => x"08",
          8690 => x"5f",
          8691 => x"ea",
          8692 => x"9c",
          8693 => x"05",
          8694 => x"5c",
          8695 => x"8d",
          8696 => x"22",
          8697 => x"b0",
          8698 => x"5d",
          8699 => x"1a",
          8700 => x"58",
          8701 => x"57",
          8702 => x"70",
          8703 => x"34",
          8704 => x"74",
          8705 => x"56",
          8706 => x"55",
          8707 => x"81",
          8708 => x"54",
          8709 => x"77",
          8710 => x"33",
          8711 => x"3f",
          8712 => x"08",
          8713 => x"81",
          8714 => x"39",
          8715 => x"0c",
          8716 => x"b8",
          8717 => x"3d",
          8718 => x"54",
          8719 => x"53",
          8720 => x"53",
          8721 => x"52",
          8722 => x"3f",
          8723 => x"08",
          8724 => x"84",
          8725 => x"83",
          8726 => x"19",
          8727 => x"08",
          8728 => x"a0",
          8729 => x"fe",
          8730 => x"19",
          8731 => x"82",
          8732 => x"06",
          8733 => x"81",
          8734 => x"08",
          8735 => x"05",
          8736 => x"81",
          8737 => x"e3",
          8738 => x"c5",
          8739 => x"22",
          8740 => x"ff",
          8741 => x"74",
          8742 => x"81",
          8743 => x"7c",
          8744 => x"fe",
          8745 => x"08",
          8746 => x"56",
          8747 => x"7d",
          8748 => x"38",
          8749 => x"76",
          8750 => x"1b",
          8751 => x"19",
          8752 => x"f8",
          8753 => x"84",
          8754 => x"8f",
          8755 => x"ee",
          8756 => x"66",
          8757 => x"7c",
          8758 => x"81",
          8759 => x"1e",
          8760 => x"5e",
          8761 => x"82",
          8762 => x"19",
          8763 => x"80",
          8764 => x"08",
          8765 => x"d1",
          8766 => x"33",
          8767 => x"74",
          8768 => x"81",
          8769 => x"38",
          8770 => x"53",
          8771 => x"81",
          8772 => x"e1",
          8773 => x"b8",
          8774 => x"2e",
          8775 => x"5a",
          8776 => x"b4",
          8777 => x"5b",
          8778 => x"38",
          8779 => x"70",
          8780 => x"76",
          8781 => x"81",
          8782 => x"33",
          8783 => x"81",
          8784 => x"41",
          8785 => x"34",
          8786 => x"32",
          8787 => x"ae",
          8788 => x"72",
          8789 => x"80",
          8790 => x"45",
          8791 => x"74",
          8792 => x"7a",
          8793 => x"56",
          8794 => x"81",
          8795 => x"60",
          8796 => x"38",
          8797 => x"80",
          8798 => x"fa",
          8799 => x"b8",
          8800 => x"84",
          8801 => x"81",
          8802 => x"1c",
          8803 => x"fe",
          8804 => x"84",
          8805 => x"94",
          8806 => x"81",
          8807 => x"08",
          8808 => x"81",
          8809 => x"e1",
          8810 => x"57",
          8811 => x"08",
          8812 => x"81",
          8813 => x"38",
          8814 => x"08",
          8815 => x"b4",
          8816 => x"1a",
          8817 => x"b8",
          8818 => x"5b",
          8819 => x"08",
          8820 => x"38",
          8821 => x"41",
          8822 => x"09",
          8823 => x"a8",
          8824 => x"b4",
          8825 => x"1a",
          8826 => x"7e",
          8827 => x"33",
          8828 => x"3f",
          8829 => x"90",
          8830 => x"2e",
          8831 => x"81",
          8832 => x"86",
          8833 => x"5b",
          8834 => x"93",
          8835 => x"33",
          8836 => x"06",
          8837 => x"08",
          8838 => x"0c",
          8839 => x"76",
          8840 => x"38",
          8841 => x"74",
          8842 => x"39",
          8843 => x"60",
          8844 => x"06",
          8845 => x"c1",
          8846 => x"80",
          8847 => x"0c",
          8848 => x"e4",
          8849 => x"0d",
          8850 => x"fd",
          8851 => x"18",
          8852 => x"77",
          8853 => x"06",
          8854 => x"19",
          8855 => x"33",
          8856 => x"71",
          8857 => x"58",
          8858 => x"ff",
          8859 => x"33",
          8860 => x"06",
          8861 => x"05",
          8862 => x"76",
          8863 => x"e4",
          8864 => x"78",
          8865 => x"33",
          8866 => x"88",
          8867 => x"44",
          8868 => x"2e",
          8869 => x"79",
          8870 => x"ff",
          8871 => x"10",
          8872 => x"5c",
          8873 => x"23",
          8874 => x"81",
          8875 => x"77",
          8876 => x"77",
          8877 => x"2a",
          8878 => x"57",
          8879 => x"90",
          8880 => x"fe",
          8881 => x"38",
          8882 => x"05",
          8883 => x"23",
          8884 => x"81",
          8885 => x"41",
          8886 => x"75",
          8887 => x"2e",
          8888 => x"ff",
          8889 => x"39",
          8890 => x"7c",
          8891 => x"74",
          8892 => x"81",
          8893 => x"78",
          8894 => x"5a",
          8895 => x"05",
          8896 => x"06",
          8897 => x"56",
          8898 => x"38",
          8899 => x"fd",
          8900 => x"0b",
          8901 => x"7a",
          8902 => x"0c",
          8903 => x"04",
          8904 => x"63",
          8905 => x"5c",
          8906 => x"51",
          8907 => x"84",
          8908 => x"5a",
          8909 => x"08",
          8910 => x"81",
          8911 => x"5d",
          8912 => x"1d",
          8913 => x"5e",
          8914 => x"56",
          8915 => x"1b",
          8916 => x"82",
          8917 => x"1b",
          8918 => x"55",
          8919 => x"09",
          8920 => x"df",
          8921 => x"75",
          8922 => x"52",
          8923 => x"51",
          8924 => x"84",
          8925 => x"80",
          8926 => x"ff",
          8927 => x"75",
          8928 => x"76",
          8929 => x"b2",
          8930 => x"08",
          8931 => x"59",
          8932 => x"84",
          8933 => x"19",
          8934 => x"70",
          8935 => x"57",
          8936 => x"1d",
          8937 => x"e5",
          8938 => x"38",
          8939 => x"81",
          8940 => x"8f",
          8941 => x"38",
          8942 => x"38",
          8943 => x"81",
          8944 => x"aa",
          8945 => x"56",
          8946 => x"74",
          8947 => x"81",
          8948 => x"78",
          8949 => x"5a",
          8950 => x"05",
          8951 => x"06",
          8952 => x"56",
          8953 => x"38",
          8954 => x"80",
          8955 => x"1c",
          8956 => x"57",
          8957 => x"8b",
          8958 => x"59",
          8959 => x"81",
          8960 => x"78",
          8961 => x"5a",
          8962 => x"31",
          8963 => x"58",
          8964 => x"80",
          8965 => x"38",
          8966 => x"e1",
          8967 => x"5d",
          8968 => x"1d",
          8969 => x"7b",
          8970 => x"3f",
          8971 => x"08",
          8972 => x"e4",
          8973 => x"fe",
          8974 => x"84",
          8975 => x"93",
          8976 => x"81",
          8977 => x"08",
          8978 => x"81",
          8979 => x"dc",
          8980 => x"57",
          8981 => x"08",
          8982 => x"81",
          8983 => x"38",
          8984 => x"08",
          8985 => x"b4",
          8986 => x"1c",
          8987 => x"b8",
          8988 => x"59",
          8989 => x"08",
          8990 => x"38",
          8991 => x"5a",
          8992 => x"09",
          8993 => x"dd",
          8994 => x"b4",
          8995 => x"1c",
          8996 => x"7d",
          8997 => x"33",
          8998 => x"3f",
          8999 => x"c5",
          9000 => x"fd",
          9001 => x"1c",
          9002 => x"2a",
          9003 => x"55",
          9004 => x"38",
          9005 => x"81",
          9006 => x"80",
          9007 => x"8d",
          9008 => x"81",
          9009 => x"90",
          9010 => x"ac",
          9011 => x"5e",
          9012 => x"2e",
          9013 => x"ff",
          9014 => x"80",
          9015 => x"f4",
          9016 => x"b8",
          9017 => x"84",
          9018 => x"80",
          9019 => x"38",
          9020 => x"75",
          9021 => x"c2",
          9022 => x"5d",
          9023 => x"1d",
          9024 => x"39",
          9025 => x"57",
          9026 => x"09",
          9027 => x"38",
          9028 => x"9b",
          9029 => x"1b",
          9030 => x"2b",
          9031 => x"40",
          9032 => x"38",
          9033 => x"bf",
          9034 => x"f3",
          9035 => x"81",
          9036 => x"83",
          9037 => x"33",
          9038 => x"11",
          9039 => x"71",
          9040 => x"52",
          9041 => x"80",
          9042 => x"38",
          9043 => x"26",
          9044 => x"76",
          9045 => x"8a",
          9046 => x"e4",
          9047 => x"61",
          9048 => x"53",
          9049 => x"5b",
          9050 => x"f6",
          9051 => x"b8",
          9052 => x"09",
          9053 => x"de",
          9054 => x"81",
          9055 => x"78",
          9056 => x"38",
          9057 => x"86",
          9058 => x"56",
          9059 => x"2e",
          9060 => x"80",
          9061 => x"79",
          9062 => x"70",
          9063 => x"7f",
          9064 => x"ff",
          9065 => x"ff",
          9066 => x"fe",
          9067 => x"0b",
          9068 => x"0c",
          9069 => x"04",
          9070 => x"ff",
          9071 => x"38",
          9072 => x"fe",
          9073 => x"3d",
          9074 => x"08",
          9075 => x"33",
          9076 => x"58",
          9077 => x"86",
          9078 => x"b5",
          9079 => x"1d",
          9080 => x"57",
          9081 => x"80",
          9082 => x"81",
          9083 => x"17",
          9084 => x"56",
          9085 => x"38",
          9086 => x"1f",
          9087 => x"60",
          9088 => x"55",
          9089 => x"05",
          9090 => x"70",
          9091 => x"34",
          9092 => x"74",
          9093 => x"80",
          9094 => x"70",
          9095 => x"56",
          9096 => x"82",
          9097 => x"c0",
          9098 => x"34",
          9099 => x"3d",
          9100 => x"1c",
          9101 => x"59",
          9102 => x"5a",
          9103 => x"70",
          9104 => x"33",
          9105 => x"05",
          9106 => x"15",
          9107 => x"38",
          9108 => x"80",
          9109 => x"79",
          9110 => x"74",
          9111 => x"38",
          9112 => x"5a",
          9113 => x"75",
          9114 => x"10",
          9115 => x"2a",
          9116 => x"ff",
          9117 => x"2a",
          9118 => x"58",
          9119 => x"80",
          9120 => x"76",
          9121 => x"32",
          9122 => x"58",
          9123 => x"d7",
          9124 => x"55",
          9125 => x"87",
          9126 => x"80",
          9127 => x"58",
          9128 => x"bf",
          9129 => x"75",
          9130 => x"87",
          9131 => x"76",
          9132 => x"ff",
          9133 => x"2a",
          9134 => x"76",
          9135 => x"1f",
          9136 => x"79",
          9137 => x"58",
          9138 => x"27",
          9139 => x"33",
          9140 => x"2e",
          9141 => x"16",
          9142 => x"27",
          9143 => x"75",
          9144 => x"56",
          9145 => x"2e",
          9146 => x"ea",
          9147 => x"56",
          9148 => x"87",
          9149 => x"98",
          9150 => x"ec",
          9151 => x"71",
          9152 => x"41",
          9153 => x"87",
          9154 => x"f4",
          9155 => x"f8",
          9156 => x"b8",
          9157 => x"38",
          9158 => x"80",
          9159 => x"fe",
          9160 => x"56",
          9161 => x"2e",
          9162 => x"84",
          9163 => x"56",
          9164 => x"08",
          9165 => x"81",
          9166 => x"38",
          9167 => x"05",
          9168 => x"34",
          9169 => x"84",
          9170 => x"05",
          9171 => x"75",
          9172 => x"06",
          9173 => x"7e",
          9174 => x"38",
          9175 => x"1d",
          9176 => x"c1",
          9177 => x"e4",
          9178 => x"80",
          9179 => x"ed",
          9180 => x"b8",
          9181 => x"84",
          9182 => x"81",
          9183 => x"b8",
          9184 => x"19",
          9185 => x"1e",
          9186 => x"57",
          9187 => x"76",
          9188 => x"38",
          9189 => x"40",
          9190 => x"09",
          9191 => x"a3",
          9192 => x"75",
          9193 => x"52",
          9194 => x"51",
          9195 => x"84",
          9196 => x"80",
          9197 => x"ff",
          9198 => x"75",
          9199 => x"76",
          9200 => x"38",
          9201 => x"70",
          9202 => x"74",
          9203 => x"81",
          9204 => x"30",
          9205 => x"78",
          9206 => x"74",
          9207 => x"c9",
          9208 => x"59",
          9209 => x"86",
          9210 => x"52",
          9211 => x"83",
          9212 => x"e4",
          9213 => x"b8",
          9214 => x"2e",
          9215 => x"87",
          9216 => x"2e",
          9217 => x"75",
          9218 => x"83",
          9219 => x"40",
          9220 => x"38",
          9221 => x"57",
          9222 => x"77",
          9223 => x"83",
          9224 => x"57",
          9225 => x"82",
          9226 => x"76",
          9227 => x"52",
          9228 => x"51",
          9229 => x"84",
          9230 => x"80",
          9231 => x"ff",
          9232 => x"76",
          9233 => x"75",
          9234 => x"c3",
          9235 => x"9c",
          9236 => x"55",
          9237 => x"81",
          9238 => x"ff",
          9239 => x"f4",
          9240 => x"9c",
          9241 => x"58",
          9242 => x"70",
          9243 => x"33",
          9244 => x"05",
          9245 => x"15",
          9246 => x"38",
          9247 => x"ab",
          9248 => x"06",
          9249 => x"8c",
          9250 => x"0b",
          9251 => x"77",
          9252 => x"b8",
          9253 => x"3d",
          9254 => x"75",
          9255 => x"25",
          9256 => x"40",
          9257 => x"b9",
          9258 => x"81",
          9259 => x"ec",
          9260 => x"b8",
          9261 => x"84",
          9262 => x"80",
          9263 => x"38",
          9264 => x"81",
          9265 => x"08",
          9266 => x"81",
          9267 => x"d3",
          9268 => x"b8",
          9269 => x"2e",
          9270 => x"83",
          9271 => x"b8",
          9272 => x"19",
          9273 => x"08",
          9274 => x"31",
          9275 => x"19",
          9276 => x"38",
          9277 => x"41",
          9278 => x"84",
          9279 => x"b8",
          9280 => x"fd",
          9281 => x"85",
          9282 => x"08",
          9283 => x"58",
          9284 => x"e9",
          9285 => x"e4",
          9286 => x"b8",
          9287 => x"ef",
          9288 => x"b8",
          9289 => x"58",
          9290 => x"81",
          9291 => x"80",
          9292 => x"70",
          9293 => x"33",
          9294 => x"70",
          9295 => x"ff",
          9296 => x"5d",
          9297 => x"74",
          9298 => x"b8",
          9299 => x"98",
          9300 => x"80",
          9301 => x"08",
          9302 => x"38",
          9303 => x"5b",
          9304 => x"09",
          9305 => x"c9",
          9306 => x"76",
          9307 => x"52",
          9308 => x"51",
          9309 => x"84",
          9310 => x"80",
          9311 => x"ff",
          9312 => x"76",
          9313 => x"75",
          9314 => x"83",
          9315 => x"08",
          9316 => x"61",
          9317 => x"5f",
          9318 => x"8d",
          9319 => x"0b",
          9320 => x"75",
          9321 => x"75",
          9322 => x"75",
          9323 => x"7c",
          9324 => x"05",
          9325 => x"58",
          9326 => x"ff",
          9327 => x"38",
          9328 => x"70",
          9329 => x"5b",
          9330 => x"e4",
          9331 => x"7b",
          9332 => x"75",
          9333 => x"57",
          9334 => x"2a",
          9335 => x"34",
          9336 => x"83",
          9337 => x"81",
          9338 => x"78",
          9339 => x"76",
          9340 => x"2e",
          9341 => x"78",
          9342 => x"22",
          9343 => x"80",
          9344 => x"38",
          9345 => x"81",
          9346 => x"34",
          9347 => x"51",
          9348 => x"84",
          9349 => x"58",
          9350 => x"08",
          9351 => x"7f",
          9352 => x"7f",
          9353 => x"fb",
          9354 => x"54",
          9355 => x"53",
          9356 => x"53",
          9357 => x"52",
          9358 => x"3f",
          9359 => x"b8",
          9360 => x"83",
          9361 => x"e4",
          9362 => x"34",
          9363 => x"a8",
          9364 => x"84",
          9365 => x"57",
          9366 => x"1d",
          9367 => x"c9",
          9368 => x"33",
          9369 => x"2e",
          9370 => x"fb",
          9371 => x"54",
          9372 => x"a0",
          9373 => x"53",
          9374 => x"1c",
          9375 => x"d1",
          9376 => x"fb",
          9377 => x"9c",
          9378 => x"33",
          9379 => x"74",
          9380 => x"09",
          9381 => x"ba",
          9382 => x"39",
          9383 => x"57",
          9384 => x"fa",
          9385 => x"d7",
          9386 => x"c0",
          9387 => x"d4",
          9388 => x"b4",
          9389 => x"61",
          9390 => x"33",
          9391 => x"3f",
          9392 => x"08",
          9393 => x"81",
          9394 => x"84",
          9395 => x"83",
          9396 => x"1c",
          9397 => x"08",
          9398 => x"a0",
          9399 => x"8a",
          9400 => x"33",
          9401 => x"2e",
          9402 => x"b8",
          9403 => x"fc",
          9404 => x"ff",
          9405 => x"7f",
          9406 => x"98",
          9407 => x"39",
          9408 => x"f7",
          9409 => x"70",
          9410 => x"80",
          9411 => x"38",
          9412 => x"81",
          9413 => x"08",
          9414 => x"05",
          9415 => x"81",
          9416 => x"ce",
          9417 => x"c1",
          9418 => x"b4",
          9419 => x"19",
          9420 => x"7c",
          9421 => x"33",
          9422 => x"3f",
          9423 => x"f3",
          9424 => x"61",
          9425 => x"5e",
          9426 => x"96",
          9427 => x"1c",
          9428 => x"82",
          9429 => x"1c",
          9430 => x"80",
          9431 => x"70",
          9432 => x"05",
          9433 => x"57",
          9434 => x"58",
          9435 => x"bc",
          9436 => x"74",
          9437 => x"81",
          9438 => x"56",
          9439 => x"38",
          9440 => x"14",
          9441 => x"ff",
          9442 => x"76",
          9443 => x"82",
          9444 => x"79",
          9445 => x"70",
          9446 => x"55",
          9447 => x"38",
          9448 => x"80",
          9449 => x"7a",
          9450 => x"5e",
          9451 => x"05",
          9452 => x"82",
          9453 => x"70",
          9454 => x"57",
          9455 => x"08",
          9456 => x"81",
          9457 => x"53",
          9458 => x"b2",
          9459 => x"2e",
          9460 => x"75",
          9461 => x"30",
          9462 => x"80",
          9463 => x"54",
          9464 => x"90",
          9465 => x"2e",
          9466 => x"77",
          9467 => x"59",
          9468 => x"58",
          9469 => x"81",
          9470 => x"81",
          9471 => x"76",
          9472 => x"38",
          9473 => x"05",
          9474 => x"81",
          9475 => x"1d",
          9476 => x"a5",
          9477 => x"f3",
          9478 => x"96",
          9479 => x"57",
          9480 => x"05",
          9481 => x"82",
          9482 => x"1c",
          9483 => x"33",
          9484 => x"89",
          9485 => x"1e",
          9486 => x"08",
          9487 => x"33",
          9488 => x"9c",
          9489 => x"11",
          9490 => x"82",
          9491 => x"90",
          9492 => x"2b",
          9493 => x"33",
          9494 => x"88",
          9495 => x"71",
          9496 => x"59",
          9497 => x"96",
          9498 => x"88",
          9499 => x"41",
          9500 => x"56",
          9501 => x"86",
          9502 => x"15",
          9503 => x"33",
          9504 => x"07",
          9505 => x"84",
          9506 => x"3d",
          9507 => x"e5",
          9508 => x"39",
          9509 => x"11",
          9510 => x"31",
          9511 => x"83",
          9512 => x"90",
          9513 => x"51",
          9514 => x"3f",
          9515 => x"08",
          9516 => x"06",
          9517 => x"75",
          9518 => x"81",
          9519 => x"b3",
          9520 => x"2a",
          9521 => x"34",
          9522 => x"34",
          9523 => x"58",
          9524 => x"1f",
          9525 => x"78",
          9526 => x"70",
          9527 => x"54",
          9528 => x"38",
          9529 => x"74",
          9530 => x"70",
          9531 => x"25",
          9532 => x"07",
          9533 => x"75",
          9534 => x"74",
          9535 => x"78",
          9536 => x"0b",
          9537 => x"56",
          9538 => x"72",
          9539 => x"33",
          9540 => x"77",
          9541 => x"88",
          9542 => x"1e",
          9543 => x"54",
          9544 => x"ff",
          9545 => x"54",
          9546 => x"a4",
          9547 => x"08",
          9548 => x"54",
          9549 => x"27",
          9550 => x"84",
          9551 => x"81",
          9552 => x"80",
          9553 => x"a0",
          9554 => x"ff",
          9555 => x"53",
          9556 => x"81",
          9557 => x"81",
          9558 => x"81",
          9559 => x"13",
          9560 => x"59",
          9561 => x"ff",
          9562 => x"b4",
          9563 => x"2a",
          9564 => x"80",
          9565 => x"80",
          9566 => x"73",
          9567 => x"5f",
          9568 => x"39",
          9569 => x"63",
          9570 => x"42",
          9571 => x"65",
          9572 => x"55",
          9573 => x"2e",
          9574 => x"53",
          9575 => x"2e",
          9576 => x"72",
          9577 => x"d9",
          9578 => x"08",
          9579 => x"73",
          9580 => x"94",
          9581 => x"55",
          9582 => x"82",
          9583 => x"42",
          9584 => x"58",
          9585 => x"70",
          9586 => x"52",
          9587 => x"73",
          9588 => x"72",
          9589 => x"ff",
          9590 => x"38",
          9591 => x"74",
          9592 => x"76",
          9593 => x"80",
          9594 => x"17",
          9595 => x"ff",
          9596 => x"af",
          9597 => x"9f",
          9598 => x"80",
          9599 => x"5b",
          9600 => x"82",
          9601 => x"80",
          9602 => x"89",
          9603 => x"ff",
          9604 => x"83",
          9605 => x"83",
          9606 => x"70",
          9607 => x"56",
          9608 => x"80",
          9609 => x"38",
          9610 => x"8f",
          9611 => x"70",
          9612 => x"ff",
          9613 => x"56",
          9614 => x"72",
          9615 => x"5b",
          9616 => x"38",
          9617 => x"26",
          9618 => x"76",
          9619 => x"74",
          9620 => x"17",
          9621 => x"81",
          9622 => x"56",
          9623 => x"80",
          9624 => x"38",
          9625 => x"81",
          9626 => x"32",
          9627 => x"80",
          9628 => x"51",
          9629 => x"72",
          9630 => x"38",
          9631 => x"46",
          9632 => x"33",
          9633 => x"af",
          9634 => x"72",
          9635 => x"70",
          9636 => x"25",
          9637 => x"54",
          9638 => x"38",
          9639 => x"0c",
          9640 => x"3d",
          9641 => x"42",
          9642 => x"26",
          9643 => x"b4",
          9644 => x"52",
          9645 => x"8d",
          9646 => x"b8",
          9647 => x"ff",
          9648 => x"73",
          9649 => x"86",
          9650 => x"b8",
          9651 => x"3d",
          9652 => x"e4",
          9653 => x"81",
          9654 => x"53",
          9655 => x"fe",
          9656 => x"39",
          9657 => x"ab",
          9658 => x"52",
          9659 => x"8d",
          9660 => x"e4",
          9661 => x"e4",
          9662 => x"0d",
          9663 => x"80",
          9664 => x"30",
          9665 => x"73",
          9666 => x"5a",
          9667 => x"2e",
          9668 => x"14",
          9669 => x"70",
          9670 => x"56",
          9671 => x"dd",
          9672 => x"dc",
          9673 => x"70",
          9674 => x"07",
          9675 => x"7d",
          9676 => x"61",
          9677 => x"27",
          9678 => x"76",
          9679 => x"f8",
          9680 => x"2e",
          9681 => x"76",
          9682 => x"80",
          9683 => x"76",
          9684 => x"fe",
          9685 => x"70",
          9686 => x"30",
          9687 => x"52",
          9688 => x"56",
          9689 => x"2e",
          9690 => x"89",
          9691 => x"57",
          9692 => x"76",
          9693 => x"56",
          9694 => x"76",
          9695 => x"c7",
          9696 => x"22",
          9697 => x"ff",
          9698 => x"5d",
          9699 => x"a0",
          9700 => x"38",
          9701 => x"ff",
          9702 => x"ae",
          9703 => x"38",
          9704 => x"aa",
          9705 => x"fe",
          9706 => x"5a",
          9707 => x"2e",
          9708 => x"10",
          9709 => x"54",
          9710 => x"76",
          9711 => x"38",
          9712 => x"22",
          9713 => x"ae",
          9714 => x"06",
          9715 => x"0b",
          9716 => x"53",
          9717 => x"81",
          9718 => x"ff",
          9719 => x"f4",
          9720 => x"5c",
          9721 => x"16",
          9722 => x"19",
          9723 => x"5d",
          9724 => x"80",
          9725 => x"a0",
          9726 => x"38",
          9727 => x"70",
          9728 => x"25",
          9729 => x"75",
          9730 => x"ce",
          9731 => x"bb",
          9732 => x"7c",
          9733 => x"38",
          9734 => x"77",
          9735 => x"70",
          9736 => x"25",
          9737 => x"51",
          9738 => x"72",
          9739 => x"e0",
          9740 => x"2e",
          9741 => x"75",
          9742 => x"38",
          9743 => x"5a",
          9744 => x"9e",
          9745 => x"88",
          9746 => x"82",
          9747 => x"06",
          9748 => x"5f",
          9749 => x"70",
          9750 => x"58",
          9751 => x"ff",
          9752 => x"1c",
          9753 => x"81",
          9754 => x"84",
          9755 => x"2e",
          9756 => x"7d",
          9757 => x"77",
          9758 => x"ed",
          9759 => x"06",
          9760 => x"2e",
          9761 => x"79",
          9762 => x"06",
          9763 => x"38",
          9764 => x"5d",
          9765 => x"85",
          9766 => x"07",
          9767 => x"2a",
          9768 => x"7d",
          9769 => x"38",
          9770 => x"5a",
          9771 => x"34",
          9772 => x"ec",
          9773 => x"e4",
          9774 => x"33",
          9775 => x"b8",
          9776 => x"2e",
          9777 => x"84",
          9778 => x"84",
          9779 => x"06",
          9780 => x"74",
          9781 => x"06",
          9782 => x"2e",
          9783 => x"74",
          9784 => x"06",
          9785 => x"98",
          9786 => x"65",
          9787 => x"42",
          9788 => x"58",
          9789 => x"ce",
          9790 => x"70",
          9791 => x"70",
          9792 => x"56",
          9793 => x"2e",
          9794 => x"80",
          9795 => x"38",
          9796 => x"5a",
          9797 => x"82",
          9798 => x"75",
          9799 => x"81",
          9800 => x"38",
          9801 => x"73",
          9802 => x"81",
          9803 => x"38",
          9804 => x"5b",
          9805 => x"80",
          9806 => x"56",
          9807 => x"76",
          9808 => x"38",
          9809 => x"75",
          9810 => x"57",
          9811 => x"53",
          9812 => x"e9",
          9813 => x"07",
          9814 => x"1d",
          9815 => x"e3",
          9816 => x"b8",
          9817 => x"1d",
          9818 => x"84",
          9819 => x"fe",
          9820 => x"82",
          9821 => x"58",
          9822 => x"38",
          9823 => x"70",
          9824 => x"06",
          9825 => x"80",
          9826 => x"38",
          9827 => x"83",
          9828 => x"05",
          9829 => x"33",
          9830 => x"33",
          9831 => x"07",
          9832 => x"57",
          9833 => x"83",
          9834 => x"38",
          9835 => x"0c",
          9836 => x"55",
          9837 => x"39",
          9838 => x"74",
          9839 => x"f0",
          9840 => x"59",
          9841 => x"38",
          9842 => x"79",
          9843 => x"17",
          9844 => x"81",
          9845 => x"2b",
          9846 => x"70",
          9847 => x"5e",
          9848 => x"09",
          9849 => x"95",
          9850 => x"07",
          9851 => x"39",
          9852 => x"1d",
          9853 => x"2e",
          9854 => x"fc",
          9855 => x"39",
          9856 => x"ab",
          9857 => x"0b",
          9858 => x"0c",
          9859 => x"04",
          9860 => x"26",
          9861 => x"ff",
          9862 => x"c9",
          9863 => x"59",
          9864 => x"81",
          9865 => x"83",
          9866 => x"18",
          9867 => x"fc",
          9868 => x"82",
          9869 => x"b5",
          9870 => x"81",
          9871 => x"84",
          9872 => x"83",
          9873 => x"70",
          9874 => x"06",
          9875 => x"80",
          9876 => x"74",
          9877 => x"83",
          9878 => x"33",
          9879 => x"81",
          9880 => x"b9",
          9881 => x"2e",
          9882 => x"83",
          9883 => x"83",
          9884 => x"70",
          9885 => x"56",
          9886 => x"80",
          9887 => x"38",
          9888 => x"8f",
          9889 => x"70",
          9890 => x"ff",
          9891 => x"59",
          9892 => x"72",
          9893 => x"59",
          9894 => x"38",
          9895 => x"54",
          9896 => x"8a",
          9897 => x"07",
          9898 => x"06",
          9899 => x"9f",
          9900 => x"99",
          9901 => x"7d",
          9902 => x"81",
          9903 => x"17",
          9904 => x"ff",
          9905 => x"5f",
          9906 => x"a0",
          9907 => x"79",
          9908 => x"5b",
          9909 => x"fa",
          9910 => x"53",
          9911 => x"83",
          9912 => x"70",
          9913 => x"5a",
          9914 => x"2e",
          9915 => x"80",
          9916 => x"07",
          9917 => x"05",
          9918 => x"74",
          9919 => x"1b",
          9920 => x"80",
          9921 => x"80",
          9922 => x"71",
          9923 => x"90",
          9924 => x"07",
          9925 => x"5a",
          9926 => x"39",
          9927 => x"05",
          9928 => x"54",
          9929 => x"34",
          9930 => x"11",
          9931 => x"5b",
          9932 => x"81",
          9933 => x"9c",
          9934 => x"07",
          9935 => x"58",
          9936 => x"e5",
          9937 => x"06",
          9938 => x"fd",
          9939 => x"82",
          9940 => x"5c",
          9941 => x"38",
          9942 => x"b8",
          9943 => x"3d",
          9944 => x"3d",
          9945 => x"02",
          9946 => x"e7",
          9947 => x"42",
          9948 => x"0c",
          9949 => x"70",
          9950 => x"79",
          9951 => x"d7",
          9952 => x"81",
          9953 => x"70",
          9954 => x"56",
          9955 => x"85",
          9956 => x"ed",
          9957 => x"2e",
          9958 => x"84",
          9959 => x"56",
          9960 => x"85",
          9961 => x"10",
          9962 => x"ac",
          9963 => x"58",
          9964 => x"76",
          9965 => x"96",
          9966 => x"0c",
          9967 => x"06",
          9968 => x"59",
          9969 => x"9b",
          9970 => x"33",
          9971 => x"b0",
          9972 => x"e4",
          9973 => x"06",
          9974 => x"5e",
          9975 => x"2e",
          9976 => x"80",
          9977 => x"16",
          9978 => x"d8",
          9979 => x"18",
          9980 => x"81",
          9981 => x"ff",
          9982 => x"84",
          9983 => x"81",
          9984 => x"81",
          9985 => x"83",
          9986 => x"c2",
          9987 => x"2e",
          9988 => x"82",
          9989 => x"41",
          9990 => x"84",
          9991 => x"5b",
          9992 => x"34",
          9993 => x"18",
          9994 => x"5a",
          9995 => x"7a",
          9996 => x"70",
          9997 => x"33",
          9998 => x"bb",
          9999 => x"b8",
         10000 => x"2e",
         10001 => x"55",
         10002 => x"b4",
         10003 => x"56",
         10004 => x"84",
         10005 => x"84",
         10006 => x"71",
         10007 => x"56",
         10008 => x"74",
         10009 => x"2e",
         10010 => x"75",
         10011 => x"38",
         10012 => x"1d",
         10013 => x"85",
         10014 => x"58",
         10015 => x"83",
         10016 => x"58",
         10017 => x"83",
         10018 => x"c4",
         10019 => x"c3",
         10020 => x"88",
         10021 => x"59",
         10022 => x"2e",
         10023 => x"83",
         10024 => x"cf",
         10025 => x"ce",
         10026 => x"88",
         10027 => x"5a",
         10028 => x"80",
         10029 => x"11",
         10030 => x"33",
         10031 => x"71",
         10032 => x"81",
         10033 => x"72",
         10034 => x"75",
         10035 => x"56",
         10036 => x"5e",
         10037 => x"a0",
         10038 => x"c8",
         10039 => x"18",
         10040 => x"17",
         10041 => x"70",
         10042 => x"5f",
         10043 => x"58",
         10044 => x"82",
         10045 => x"81",
         10046 => x"71",
         10047 => x"19",
         10048 => x"5a",
         10049 => x"23",
         10050 => x"80",
         10051 => x"38",
         10052 => x"06",
         10053 => x"bb",
         10054 => x"17",
         10055 => x"18",
         10056 => x"2b",
         10057 => x"74",
         10058 => x"74",
         10059 => x"5e",
         10060 => x"7c",
         10061 => x"80",
         10062 => x"80",
         10063 => x"71",
         10064 => x"56",
         10065 => x"38",
         10066 => x"83",
         10067 => x"12",
         10068 => x"2b",
         10069 => x"07",
         10070 => x"70",
         10071 => x"2b",
         10072 => x"07",
         10073 => x"58",
         10074 => x"80",
         10075 => x"80",
         10076 => x"71",
         10077 => x"5d",
         10078 => x"7b",
         10079 => x"ce",
         10080 => x"7a",
         10081 => x"5a",
         10082 => x"81",
         10083 => x"52",
         10084 => x"51",
         10085 => x"3f",
         10086 => x"08",
         10087 => x"e4",
         10088 => x"81",
         10089 => x"b8",
         10090 => x"ff",
         10091 => x"26",
         10092 => x"5d",
         10093 => x"f5",
         10094 => x"82",
         10095 => x"f5",
         10096 => x"38",
         10097 => x"16",
         10098 => x"0c",
         10099 => x"0c",
         10100 => x"a8",
         10101 => x"1d",
         10102 => x"57",
         10103 => x"2e",
         10104 => x"88",
         10105 => x"8d",
         10106 => x"2e",
         10107 => x"7d",
         10108 => x"0c",
         10109 => x"7c",
         10110 => x"38",
         10111 => x"70",
         10112 => x"81",
         10113 => x"5a",
         10114 => x"89",
         10115 => x"58",
         10116 => x"08",
         10117 => x"ff",
         10118 => x"0c",
         10119 => x"18",
         10120 => x"0b",
         10121 => x"7c",
         10122 => x"96",
         10123 => x"34",
         10124 => x"22",
         10125 => x"7c",
         10126 => x"23",
         10127 => x"23",
         10128 => x"0b",
         10129 => x"80",
         10130 => x"0c",
         10131 => x"84",
         10132 => x"97",
         10133 => x"8b",
         10134 => x"e4",
         10135 => x"0d",
         10136 => x"d0",
         10137 => x"ff",
         10138 => x"58",
         10139 => x"91",
         10140 => x"78",
         10141 => x"d0",
         10142 => x"78",
         10143 => x"fe",
         10144 => x"08",
         10145 => x"5f",
         10146 => x"08",
         10147 => x"7a",
         10148 => x"5c",
         10149 => x"81",
         10150 => x"ff",
         10151 => x"58",
         10152 => x"26",
         10153 => x"16",
         10154 => x"06",
         10155 => x"9f",
         10156 => x"99",
         10157 => x"e0",
         10158 => x"ff",
         10159 => x"75",
         10160 => x"2a",
         10161 => x"77",
         10162 => x"06",
         10163 => x"ff",
         10164 => x"7a",
         10165 => x"70",
         10166 => x"2a",
         10167 => x"58",
         10168 => x"2e",
         10169 => x"81",
         10170 => x"5e",
         10171 => x"25",
         10172 => x"61",
         10173 => x"39",
         10174 => x"fe",
         10175 => x"82",
         10176 => x"5e",
         10177 => x"fe",
         10178 => x"58",
         10179 => x"7a",
         10180 => x"59",
         10181 => x"2e",
         10182 => x"83",
         10183 => x"75",
         10184 => x"70",
         10185 => x"25",
         10186 => x"5b",
         10187 => x"ad",
         10188 => x"e8",
         10189 => x"38",
         10190 => x"57",
         10191 => x"83",
         10192 => x"70",
         10193 => x"80",
         10194 => x"84",
         10195 => x"84",
         10196 => x"71",
         10197 => x"88",
         10198 => x"ff",
         10199 => x"72",
         10200 => x"83",
         10201 => x"71",
         10202 => x"5b",
         10203 => x"77",
         10204 => x"05",
         10205 => x"19",
         10206 => x"59",
         10207 => x"ff",
         10208 => x"b8",
         10209 => x"70",
         10210 => x"2a",
         10211 => x"9b",
         10212 => x"10",
         10213 => x"84",
         10214 => x"5d",
         10215 => x"42",
         10216 => x"83",
         10217 => x"2e",
         10218 => x"80",
         10219 => x"34",
         10220 => x"18",
         10221 => x"80",
         10222 => x"2e",
         10223 => x"54",
         10224 => x"17",
         10225 => x"33",
         10226 => x"86",
         10227 => x"e4",
         10228 => x"85",
         10229 => x"81",
         10230 => x"18",
         10231 => x"75",
         10232 => x"1f",
         10233 => x"71",
         10234 => x"5d",
         10235 => x"7b",
         10236 => x"2e",
         10237 => x"a8",
         10238 => x"b8",
         10239 => x"58",
         10240 => x"2e",
         10241 => x"75",
         10242 => x"70",
         10243 => x"25",
         10244 => x"42",
         10245 => x"38",
         10246 => x"2e",
         10247 => x"58",
         10248 => x"06",
         10249 => x"84",
         10250 => x"33",
         10251 => x"78",
         10252 => x"06",
         10253 => x"58",
         10254 => x"f8",
         10255 => x"80",
         10256 => x"38",
         10257 => x"1a",
         10258 => x"7a",
         10259 => x"38",
         10260 => x"83",
         10261 => x"18",
         10262 => x"40",
         10263 => x"70",
         10264 => x"33",
         10265 => x"05",
         10266 => x"71",
         10267 => x"5b",
         10268 => x"77",
         10269 => x"c5",
         10270 => x"2e",
         10271 => x"0b",
         10272 => x"83",
         10273 => x"5d",
         10274 => x"81",
         10275 => x"7e",
         10276 => x"40",
         10277 => x"31",
         10278 => x"58",
         10279 => x"80",
         10280 => x"38",
         10281 => x"e1",
         10282 => x"fe",
         10283 => x"58",
         10284 => x"38",
         10285 => x"e4",
         10286 => x"0d",
         10287 => x"75",
         10288 => x"dc",
         10289 => x"81",
         10290 => x"e4",
         10291 => x"58",
         10292 => x"8d",
         10293 => x"e4",
         10294 => x"0d",
         10295 => x"80",
         10296 => x"e4",
         10297 => x"58",
         10298 => x"05",
         10299 => x"70",
         10300 => x"33",
         10301 => x"ff",
         10302 => x"5f",
         10303 => x"2e",
         10304 => x"74",
         10305 => x"38",
         10306 => x"8a",
         10307 => x"98",
         10308 => x"78",
         10309 => x"5a",
         10310 => x"81",
         10311 => x"71",
         10312 => x"1b",
         10313 => x"40",
         10314 => x"84",
         10315 => x"80",
         10316 => x"93",
         10317 => x"5a",
         10318 => x"83",
         10319 => x"fd",
         10320 => x"e9",
         10321 => x"e8",
         10322 => x"88",
         10323 => x"55",
         10324 => x"09",
         10325 => x"d5",
         10326 => x"58",
         10327 => x"17",
         10328 => x"b1",
         10329 => x"33",
         10330 => x"2e",
         10331 => x"82",
         10332 => x"54",
         10333 => x"17",
         10334 => x"33",
         10335 => x"d2",
         10336 => x"e4",
         10337 => x"85",
         10338 => x"81",
         10339 => x"18",
         10340 => x"99",
         10341 => x"18",
         10342 => x"17",
         10343 => x"18",
         10344 => x"2b",
         10345 => x"75",
         10346 => x"2e",
         10347 => x"f8",
         10348 => x"17",
         10349 => x"82",
         10350 => x"90",
         10351 => x"2b",
         10352 => x"33",
         10353 => x"88",
         10354 => x"71",
         10355 => x"59",
         10356 => x"59",
         10357 => x"85",
         10358 => x"09",
         10359 => x"cd",
         10360 => x"17",
         10361 => x"82",
         10362 => x"90",
         10363 => x"2b",
         10364 => x"33",
         10365 => x"88",
         10366 => x"71",
         10367 => x"40",
         10368 => x"5e",
         10369 => x"85",
         10370 => x"09",
         10371 => x"9d",
         10372 => x"17",
         10373 => x"82",
         10374 => x"90",
         10375 => x"2b",
         10376 => x"33",
         10377 => x"88",
         10378 => x"71",
         10379 => x"0c",
         10380 => x"1c",
         10381 => x"82",
         10382 => x"90",
         10383 => x"2b",
         10384 => x"33",
         10385 => x"88",
         10386 => x"71",
         10387 => x"05",
         10388 => x"49",
         10389 => x"40",
         10390 => x"5a",
         10391 => x"84",
         10392 => x"81",
         10393 => x"84",
         10394 => x"7c",
         10395 => x"84",
         10396 => x"8c",
         10397 => x"0b",
         10398 => x"f7",
         10399 => x"83",
         10400 => x"38",
         10401 => x"0c",
         10402 => x"39",
         10403 => x"17",
         10404 => x"17",
         10405 => x"18",
         10406 => x"ff",
         10407 => x"84",
         10408 => x"7a",
         10409 => x"06",
         10410 => x"84",
         10411 => x"83",
         10412 => x"17",
         10413 => x"08",
         10414 => x"a0",
         10415 => x"8b",
         10416 => x"33",
         10417 => x"2e",
         10418 => x"84",
         10419 => x"5a",
         10420 => x"74",
         10421 => x"2e",
         10422 => x"85",
         10423 => x"18",
         10424 => x"5c",
         10425 => x"ab",
         10426 => x"17",
         10427 => x"18",
         10428 => x"2b",
         10429 => x"8d",
         10430 => x"d2",
         10431 => x"22",
         10432 => x"ca",
         10433 => x"17",
         10434 => x"82",
         10435 => x"90",
         10436 => x"2b",
         10437 => x"33",
         10438 => x"88",
         10439 => x"71",
         10440 => x"0c",
         10441 => x"2b",
         10442 => x"40",
         10443 => x"d8",
         10444 => x"75",
         10445 => x"e8",
         10446 => x"f9",
         10447 => x"80",
         10448 => x"38",
         10449 => x"57",
         10450 => x"f7",
         10451 => x"5a",
         10452 => x"38",
         10453 => x"75",
         10454 => x"08",
         10455 => x"05",
         10456 => x"81",
         10457 => x"ff",
         10458 => x"fc",
         10459 => x"3d",
         10460 => x"d3",
         10461 => x"70",
         10462 => x"41",
         10463 => x"76",
         10464 => x"80",
         10465 => x"38",
         10466 => x"05",
         10467 => x"9f",
         10468 => x"74",
         10469 => x"e2",
         10470 => x"38",
         10471 => x"80",
         10472 => x"d0",
         10473 => x"80",
         10474 => x"c4",
         10475 => x"10",
         10476 => x"05",
         10477 => x"55",
         10478 => x"84",
         10479 => x"34",
         10480 => x"80",
         10481 => x"80",
         10482 => x"54",
         10483 => x"7c",
         10484 => x"2e",
         10485 => x"53",
         10486 => x"53",
         10487 => x"ef",
         10488 => x"b8",
         10489 => x"73",
         10490 => x"0c",
         10491 => x"04",
         10492 => x"b8",
         10493 => x"3d",
         10494 => x"33",
         10495 => x"81",
         10496 => x"56",
         10497 => x"26",
         10498 => x"16",
         10499 => x"06",
         10500 => x"58",
         10501 => x"80",
         10502 => x"7f",
         10503 => x"d4",
         10504 => x"7b",
         10505 => x"5a",
         10506 => x"05",
         10507 => x"70",
         10508 => x"33",
         10509 => x"59",
         10510 => x"99",
         10511 => x"e0",
         10512 => x"ff",
         10513 => x"ff",
         10514 => x"76",
         10515 => x"38",
         10516 => x"81",
         10517 => x"54",
         10518 => x"9f",
         10519 => x"74",
         10520 => x"81",
         10521 => x"76",
         10522 => x"77",
         10523 => x"30",
         10524 => x"9f",
         10525 => x"5c",
         10526 => x"80",
         10527 => x"81",
         10528 => x"5d",
         10529 => x"25",
         10530 => x"7f",
         10531 => x"39",
         10532 => x"f7",
         10533 => x"60",
         10534 => x"8b",
         10535 => x"0d",
         10536 => x"05",
         10537 => x"33",
         10538 => x"56",
         10539 => x"a6",
         10540 => x"06",
         10541 => x"3d",
         10542 => x"9e",
         10543 => x"52",
         10544 => x"3f",
         10545 => x"08",
         10546 => x"e4",
         10547 => x"8f",
         10548 => x"0c",
         10549 => x"84",
         10550 => x"9c",
         10551 => x"7e",
         10552 => x"90",
         10553 => x"5a",
         10554 => x"84",
         10555 => x"57",
         10556 => x"08",
         10557 => x"ba",
         10558 => x"06",
         10559 => x"2e",
         10560 => x"76",
         10561 => x"c1",
         10562 => x"2e",
         10563 => x"77",
         10564 => x"76",
         10565 => x"77",
         10566 => x"06",
         10567 => x"2e",
         10568 => x"66",
         10569 => x"9a",
         10570 => x"88",
         10571 => x"70",
         10572 => x"5e",
         10573 => x"83",
         10574 => x"38",
         10575 => x"17",
         10576 => x"8f",
         10577 => x"0b",
         10578 => x"80",
         10579 => x"17",
         10580 => x"a0",
         10581 => x"34",
         10582 => x"5e",
         10583 => x"17",
         10584 => x"9b",
         10585 => x"33",
         10586 => x"2e",
         10587 => x"66",
         10588 => x"9c",
         10589 => x"0b",
         10590 => x"80",
         10591 => x"34",
         10592 => x"1c",
         10593 => x"81",
         10594 => x"34",
         10595 => x"80",
         10596 => x"b4",
         10597 => x"7c",
         10598 => x"5f",
         10599 => x"27",
         10600 => x"17",
         10601 => x"83",
         10602 => x"57",
         10603 => x"fe",
         10604 => x"80",
         10605 => x"70",
         10606 => x"5b",
         10607 => x"fe",
         10608 => x"78",
         10609 => x"57",
         10610 => x"38",
         10611 => x"38",
         10612 => x"05",
         10613 => x"2a",
         10614 => x"56",
         10615 => x"38",
         10616 => x"81",
         10617 => x"80",
         10618 => x"75",
         10619 => x"79",
         10620 => x"77",
         10621 => x"06",
         10622 => x"2e",
         10623 => x"80",
         10624 => x"7e",
         10625 => x"a0",
         10626 => x"a4",
         10627 => x"9b",
         10628 => x"12",
         10629 => x"2b",
         10630 => x"40",
         10631 => x"5a",
         10632 => x"81",
         10633 => x"88",
         10634 => x"16",
         10635 => x"82",
         10636 => x"90",
         10637 => x"2b",
         10638 => x"33",
         10639 => x"88",
         10640 => x"71",
         10641 => x"8c",
         10642 => x"60",
         10643 => x"41",
         10644 => x"5e",
         10645 => x"84",
         10646 => x"90",
         10647 => x"0b",
         10648 => x"80",
         10649 => x"0c",
         10650 => x"81",
         10651 => x"80",
         10652 => x"38",
         10653 => x"84",
         10654 => x"94",
         10655 => x"1a",
         10656 => x"2b",
         10657 => x"58",
         10658 => x"78",
         10659 => x"56",
         10660 => x"27",
         10661 => x"81",
         10662 => x"5f",
         10663 => x"2e",
         10664 => x"77",
         10665 => x"ff",
         10666 => x"84",
         10667 => x"58",
         10668 => x"08",
         10669 => x"38",
         10670 => x"b8",
         10671 => x"2e",
         10672 => x"75",
         10673 => x"c0",
         10674 => x"c2",
         10675 => x"06",
         10676 => x"38",
         10677 => x"81",
         10678 => x"80",
         10679 => x"38",
         10680 => x"79",
         10681 => x"39",
         10682 => x"79",
         10683 => x"39",
         10684 => x"79",
         10685 => x"39",
         10686 => x"ca",
         10687 => x"e4",
         10688 => x"07",
         10689 => x"fb",
         10690 => x"8b",
         10691 => x"7b",
         10692 => x"fe",
         10693 => x"16",
         10694 => x"33",
         10695 => x"71",
         10696 => x"7d",
         10697 => x"5c",
         10698 => x"7c",
         10699 => x"27",
         10700 => x"74",
         10701 => x"ff",
         10702 => x"84",
         10703 => x"5d",
         10704 => x"08",
         10705 => x"a7",
         10706 => x"e4",
         10707 => x"fc",
         10708 => x"b8",
         10709 => x"2e",
         10710 => x"80",
         10711 => x"76",
         10712 => x"82",
         10713 => x"e4",
         10714 => x"38",
         10715 => x"fe",
         10716 => x"08",
         10717 => x"75",
         10718 => x"af",
         10719 => x"94",
         10720 => x"17",
         10721 => x"55",
         10722 => x"34",
         10723 => x"7d",
         10724 => x"38",
         10725 => x"80",
         10726 => x"34",
         10727 => x"17",
         10728 => x"39",
         10729 => x"94",
         10730 => x"98",
         10731 => x"2b",
         10732 => x"5e",
         10733 => x"0b",
         10734 => x"80",
         10735 => x"34",
         10736 => x"17",
         10737 => x"0b",
         10738 => x"66",
         10739 => x"8b",
         10740 => x"67",
         10741 => x"0b",
         10742 => x"80",
         10743 => x"34",
         10744 => x"7c",
         10745 => x"81",
         10746 => x"38",
         10747 => x"80",
         10748 => x"5e",
         10749 => x"b4",
         10750 => x"2e",
         10751 => x"16",
         10752 => x"7d",
         10753 => x"06",
         10754 => x"54",
         10755 => x"16",
         10756 => x"33",
         10757 => x"ba",
         10758 => x"e4",
         10759 => x"85",
         10760 => x"81",
         10761 => x"17",
         10762 => x"7a",
         10763 => x"18",
         10764 => x"80",
         10765 => x"38",
         10766 => x"f9",
         10767 => x"54",
         10768 => x"53",
         10769 => x"53",
         10770 => x"52",
         10771 => x"81",
         10772 => x"e4",
         10773 => x"09",
         10774 => x"aa",
         10775 => x"e4",
         10776 => x"34",
         10777 => x"a8",
         10778 => x"84",
         10779 => x"5c",
         10780 => x"17",
         10781 => x"92",
         10782 => x"33",
         10783 => x"2e",
         10784 => x"ff",
         10785 => x"54",
         10786 => x"a0",
         10787 => x"53",
         10788 => x"16",
         10789 => x"a3",
         10790 => x"5b",
         10791 => x"74",
         10792 => x"76",
         10793 => x"39",
         10794 => x"0c",
         10795 => x"38",
         10796 => x"06",
         10797 => x"2e",
         10798 => x"7e",
         10799 => x"12",
         10800 => x"5f",
         10801 => x"7d",
         10802 => x"38",
         10803 => x"78",
         10804 => x"1c",
         10805 => x"5c",
         10806 => x"f9",
         10807 => x"89",
         10808 => x"1a",
         10809 => x"f7",
         10810 => x"94",
         10811 => x"56",
         10812 => x"81",
         10813 => x"0c",
         10814 => x"84",
         10815 => x"57",
         10816 => x"f7",
         10817 => x"7f",
         10818 => x"9f",
         10819 => x"0d",
         10820 => x"66",
         10821 => x"5a",
         10822 => x"89",
         10823 => x"2e",
         10824 => x"08",
         10825 => x"2e",
         10826 => x"33",
         10827 => x"2e",
         10828 => x"16",
         10829 => x"22",
         10830 => x"78",
         10831 => x"38",
         10832 => x"41",
         10833 => x"82",
         10834 => x"1a",
         10835 => x"82",
         10836 => x"1a",
         10837 => x"57",
         10838 => x"80",
         10839 => x"38",
         10840 => x"8c",
         10841 => x"31",
         10842 => x"75",
         10843 => x"38",
         10844 => x"81",
         10845 => x"59",
         10846 => x"06",
         10847 => x"e3",
         10848 => x"22",
         10849 => x"89",
         10850 => x"7a",
         10851 => x"83",
         10852 => x"1a",
         10853 => x"75",
         10854 => x"38",
         10855 => x"83",
         10856 => x"98",
         10857 => x"59",
         10858 => x"fe",
         10859 => x"08",
         10860 => x"57",
         10861 => x"83",
         10862 => x"19",
         10863 => x"29",
         10864 => x"05",
         10865 => x"80",
         10866 => x"38",
         10867 => x"89",
         10868 => x"77",
         10869 => x"81",
         10870 => x"55",
         10871 => x"85",
         10872 => x"31",
         10873 => x"76",
         10874 => x"81",
         10875 => x"ff",
         10876 => x"84",
         10877 => x"83",
         10878 => x"83",
         10879 => x"59",
         10880 => x"a9",
         10881 => x"08",
         10882 => x"75",
         10883 => x"38",
         10884 => x"71",
         10885 => x"1b",
         10886 => x"75",
         10887 => x"57",
         10888 => x"81",
         10889 => x"ff",
         10890 => x"ef",
         10891 => x"2b",
         10892 => x"31",
         10893 => x"7f",
         10894 => x"94",
         10895 => x"70",
         10896 => x"0c",
         10897 => x"fe",
         10898 => x"56",
         10899 => x"e4",
         10900 => x"0d",
         10901 => x"b8",
         10902 => x"3d",
         10903 => x"5c",
         10904 => x"9c",
         10905 => x"75",
         10906 => x"84",
         10907 => x"59",
         10908 => x"27",
         10909 => x"58",
         10910 => x"19",
         10911 => x"b6",
         10912 => x"83",
         10913 => x"5d",
         10914 => x"7f",
         10915 => x"06",
         10916 => x"81",
         10917 => x"b8",
         10918 => x"19",
         10919 => x"9e",
         10920 => x"b8",
         10921 => x"2e",
         10922 => x"56",
         10923 => x"b4",
         10924 => x"81",
         10925 => x"94",
         10926 => x"ff",
         10927 => x"7f",
         10928 => x"05",
         10929 => x"80",
         10930 => x"38",
         10931 => x"05",
         10932 => x"70",
         10933 => x"34",
         10934 => x"75",
         10935 => x"d1",
         10936 => x"81",
         10937 => x"77",
         10938 => x"59",
         10939 => x"56",
         10940 => x"fe",
         10941 => x"54",
         10942 => x"53",
         10943 => x"53",
         10944 => x"52",
         10945 => x"c9",
         10946 => x"84",
         10947 => x"7f",
         10948 => x"06",
         10949 => x"84",
         10950 => x"83",
         10951 => x"19",
         10952 => x"08",
         10953 => x"e4",
         10954 => x"74",
         10955 => x"27",
         10956 => x"82",
         10957 => x"74",
         10958 => x"81",
         10959 => x"38",
         10960 => x"19",
         10961 => x"08",
         10962 => x"52",
         10963 => x"51",
         10964 => x"3f",
         10965 => x"bb",
         10966 => x"1b",
         10967 => x"08",
         10968 => x"39",
         10969 => x"52",
         10970 => x"a3",
         10971 => x"b8",
         10972 => x"fc",
         10973 => x"16",
         10974 => x"9c",
         10975 => x"b8",
         10976 => x"06",
         10977 => x"b8",
         10978 => x"08",
         10979 => x"b2",
         10980 => x"91",
         10981 => x"0b",
         10982 => x"0c",
         10983 => x"04",
         10984 => x"1b",
         10985 => x"84",
         10986 => x"92",
         10987 => x"f0",
         10988 => x"65",
         10989 => x"40",
         10990 => x"7e",
         10991 => x"79",
         10992 => x"38",
         10993 => x"75",
         10994 => x"38",
         10995 => x"74",
         10996 => x"38",
         10997 => x"84",
         10998 => x"59",
         10999 => x"85",
         11000 => x"55",
         11001 => x"55",
         11002 => x"38",
         11003 => x"55",
         11004 => x"38",
         11005 => x"70",
         11006 => x"06",
         11007 => x"56",
         11008 => x"82",
         11009 => x"1a",
         11010 => x"5d",
         11011 => x"27",
         11012 => x"09",
         11013 => x"2e",
         11014 => x"76",
         11015 => x"5f",
         11016 => x"38",
         11017 => x"22",
         11018 => x"89",
         11019 => x"56",
         11020 => x"76",
         11021 => x"88",
         11022 => x"74",
         11023 => x"b1",
         11024 => x"2e",
         11025 => x"74",
         11026 => x"8c",
         11027 => x"1b",
         11028 => x"08",
         11029 => x"88",
         11030 => x"56",
         11031 => x"9c",
         11032 => x"81",
         11033 => x"1a",
         11034 => x"9c",
         11035 => x"05",
         11036 => x"77",
         11037 => x"38",
         11038 => x"70",
         11039 => x"18",
         11040 => x"57",
         11041 => x"85",
         11042 => x"15",
         11043 => x"59",
         11044 => x"2e",
         11045 => x"77",
         11046 => x"7f",
         11047 => x"76",
         11048 => x"77",
         11049 => x"7c",
         11050 => x"33",
         11051 => x"a1",
         11052 => x"e4",
         11053 => x"38",
         11054 => x"08",
         11055 => x"57",
         11056 => x"a5",
         11057 => x"0b",
         11058 => x"72",
         11059 => x"58",
         11060 => x"81",
         11061 => x"77",
         11062 => x"59",
         11063 => x"56",
         11064 => x"60",
         11065 => x"1a",
         11066 => x"2b",
         11067 => x"31",
         11068 => x"7f",
         11069 => x"94",
         11070 => x"70",
         11071 => x"0c",
         11072 => x"5a",
         11073 => x"5b",
         11074 => x"83",
         11075 => x"75",
         11076 => x"7a",
         11077 => x"90",
         11078 => x"77",
         11079 => x"5b",
         11080 => x"34",
         11081 => x"84",
         11082 => x"92",
         11083 => x"74",
         11084 => x"0c",
         11085 => x"04",
         11086 => x"55",
         11087 => x"38",
         11088 => x"a2",
         11089 => x"1b",
         11090 => x"76",
         11091 => x"84",
         11092 => x"5a",
         11093 => x"27",
         11094 => x"59",
         11095 => x"16",
         11096 => x"b6",
         11097 => x"83",
         11098 => x"5e",
         11099 => x"7f",
         11100 => x"06",
         11101 => x"81",
         11102 => x"b8",
         11103 => x"16",
         11104 => x"98",
         11105 => x"b8",
         11106 => x"2e",
         11107 => x"57",
         11108 => x"b4",
         11109 => x"83",
         11110 => x"94",
         11111 => x"ff",
         11112 => x"58",
         11113 => x"59",
         11114 => x"80",
         11115 => x"76",
         11116 => x"58",
         11117 => x"81",
         11118 => x"ff",
         11119 => x"ef",
         11120 => x"81",
         11121 => x"34",
         11122 => x"81",
         11123 => x"08",
         11124 => x"70",
         11125 => x"33",
         11126 => x"98",
         11127 => x"5c",
         11128 => x"08",
         11129 => x"81",
         11130 => x"38",
         11131 => x"08",
         11132 => x"b4",
         11133 => x"17",
         11134 => x"b8",
         11135 => x"55",
         11136 => x"08",
         11137 => x"38",
         11138 => x"55",
         11139 => x"09",
         11140 => x"e3",
         11141 => x"b4",
         11142 => x"17",
         11143 => x"7f",
         11144 => x"33",
         11145 => x"a9",
         11146 => x"fe",
         11147 => x"1a",
         11148 => x"1a",
         11149 => x"93",
         11150 => x"33",
         11151 => x"b9",
         11152 => x"b4",
         11153 => x"1b",
         11154 => x"7b",
         11155 => x"0c",
         11156 => x"39",
         11157 => x"52",
         11158 => x"ab",
         11159 => x"b8",
         11160 => x"84",
         11161 => x"fb",
         11162 => x"1a",
         11163 => x"ab",
         11164 => x"79",
         11165 => x"cc",
         11166 => x"e4",
         11167 => x"b8",
         11168 => x"bd",
         11169 => x"81",
         11170 => x"08",
         11171 => x"70",
         11172 => x"33",
         11173 => x"97",
         11174 => x"b8",
         11175 => x"b8",
         11176 => x"e4",
         11177 => x"34",
         11178 => x"a8",
         11179 => x"58",
         11180 => x"08",
         11181 => x"38",
         11182 => x"5c",
         11183 => x"09",
         11184 => x"fc",
         11185 => x"b4",
         11186 => x"17",
         11187 => x"76",
         11188 => x"33",
         11189 => x"f9",
         11190 => x"fb",
         11191 => x"16",
         11192 => x"95",
         11193 => x"b8",
         11194 => x"06",
         11195 => x"f2",
         11196 => x"08",
         11197 => x"ec",
         11198 => x"b4",
         11199 => x"b8",
         11200 => x"81",
         11201 => x"57",
         11202 => x"3f",
         11203 => x"08",
         11204 => x"84",
         11205 => x"83",
         11206 => x"16",
         11207 => x"08",
         11208 => x"a0",
         11209 => x"fe",
         11210 => x"16",
         11211 => x"82",
         11212 => x"06",
         11213 => x"81",
         11214 => x"08",
         11215 => x"05",
         11216 => x"81",
         11217 => x"ff",
         11218 => x"60",
         11219 => x"0c",
         11220 => x"58",
         11221 => x"39",
         11222 => x"1b",
         11223 => x"84",
         11224 => x"92",
         11225 => x"82",
         11226 => x"34",
         11227 => x"b8",
         11228 => x"3d",
         11229 => x"3d",
         11230 => x"89",
         11231 => x"2e",
         11232 => x"08",
         11233 => x"2e",
         11234 => x"33",
         11235 => x"2e",
         11236 => x"16",
         11237 => x"22",
         11238 => x"77",
         11239 => x"38",
         11240 => x"5c",
         11241 => x"81",
         11242 => x"18",
         11243 => x"2a",
         11244 => x"57",
         11245 => x"81",
         11246 => x"a0",
         11247 => x"57",
         11248 => x"79",
         11249 => x"83",
         11250 => x"7a",
         11251 => x"81",
         11252 => x"b8",
         11253 => x"17",
         11254 => x"93",
         11255 => x"b8",
         11256 => x"2e",
         11257 => x"59",
         11258 => x"b4",
         11259 => x"81",
         11260 => x"18",
         11261 => x"33",
         11262 => x"57",
         11263 => x"34",
         11264 => x"19",
         11265 => x"ff",
         11266 => x"5a",
         11267 => x"18",
         11268 => x"2a",
         11269 => x"18",
         11270 => x"76",
         11271 => x"5c",
         11272 => x"83",
         11273 => x"38",
         11274 => x"55",
         11275 => x"74",
         11276 => x"7a",
         11277 => x"74",
         11278 => x"75",
         11279 => x"74",
         11280 => x"78",
         11281 => x"80",
         11282 => x"0b",
         11283 => x"a1",
         11284 => x"34",
         11285 => x"99",
         11286 => x"0b",
         11287 => x"80",
         11288 => x"34",
         11289 => x"0b",
         11290 => x"7b",
         11291 => x"94",
         11292 => x"e4",
         11293 => x"33",
         11294 => x"5b",
         11295 => x"19",
         11296 => x"b8",
         11297 => x"3d",
         11298 => x"54",
         11299 => x"53",
         11300 => x"53",
         11301 => x"52",
         11302 => x"b5",
         11303 => x"84",
         11304 => x"fe",
         11305 => x"b8",
         11306 => x"18",
         11307 => x"08",
         11308 => x"31",
         11309 => x"08",
         11310 => x"a0",
         11311 => x"fe",
         11312 => x"17",
         11313 => x"82",
         11314 => x"06",
         11315 => x"81",
         11316 => x"08",
         11317 => x"05",
         11318 => x"81",
         11319 => x"ff",
         11320 => x"79",
         11321 => x"39",
         11322 => x"55",
         11323 => x"34",
         11324 => x"56",
         11325 => x"34",
         11326 => x"55",
         11327 => x"74",
         11328 => x"7a",
         11329 => x"74",
         11330 => x"75",
         11331 => x"74",
         11332 => x"78",
         11333 => x"80",
         11334 => x"0b",
         11335 => x"a1",
         11336 => x"34",
         11337 => x"99",
         11338 => x"0b",
         11339 => x"80",
         11340 => x"34",
         11341 => x"0b",
         11342 => x"7b",
         11343 => x"c4",
         11344 => x"e4",
         11345 => x"33",
         11346 => x"5b",
         11347 => x"19",
         11348 => x"39",
         11349 => x"51",
         11350 => x"3f",
         11351 => x"08",
         11352 => x"74",
         11353 => x"74",
         11354 => x"5a",
         11355 => x"f9",
         11356 => x"70",
         11357 => x"fe",
         11358 => x"e4",
         11359 => x"b8",
         11360 => x"38",
         11361 => x"80",
         11362 => x"74",
         11363 => x"80",
         11364 => x"72",
         11365 => x"80",
         11366 => x"86",
         11367 => x"16",
         11368 => x"71",
         11369 => x"38",
         11370 => x"58",
         11371 => x"84",
         11372 => x"0c",
         11373 => x"e4",
         11374 => x"0d",
         11375 => x"33",
         11376 => x"bc",
         11377 => x"e4",
         11378 => x"53",
         11379 => x"73",
         11380 => x"56",
         11381 => x"3d",
         11382 => x"70",
         11383 => x"75",
         11384 => x"38",
         11385 => x"05",
         11386 => x"9f",
         11387 => x"71",
         11388 => x"38",
         11389 => x"71",
         11390 => x"38",
         11391 => x"33",
         11392 => x"24",
         11393 => x"84",
         11394 => x"80",
         11395 => x"e4",
         11396 => x"0d",
         11397 => x"84",
         11398 => x"8c",
         11399 => x"78",
         11400 => x"70",
         11401 => x"53",
         11402 => x"89",
         11403 => x"82",
         11404 => x"ff",
         11405 => x"59",
         11406 => x"2e",
         11407 => x"80",
         11408 => x"d4",
         11409 => x"08",
         11410 => x"76",
         11411 => x"58",
         11412 => x"81",
         11413 => x"ff",
         11414 => x"54",
         11415 => x"26",
         11416 => x"12",
         11417 => x"06",
         11418 => x"9f",
         11419 => x"99",
         11420 => x"e0",
         11421 => x"ff",
         11422 => x"71",
         11423 => x"2a",
         11424 => x"73",
         11425 => x"06",
         11426 => x"ff",
         11427 => x"76",
         11428 => x"70",
         11429 => x"2a",
         11430 => x"52",
         11431 => x"2e",
         11432 => x"18",
         11433 => x"58",
         11434 => x"ff",
         11435 => x"51",
         11436 => x"77",
         11437 => x"38",
         11438 => x"51",
         11439 => x"ea",
         11440 => x"53",
         11441 => x"05",
         11442 => x"51",
         11443 => x"84",
         11444 => x"55",
         11445 => x"08",
         11446 => x"38",
         11447 => x"e4",
         11448 => x"0d",
         11449 => x"68",
         11450 => x"d0",
         11451 => x"94",
         11452 => x"e4",
         11453 => x"b8",
         11454 => x"c6",
         11455 => x"d7",
         11456 => x"98",
         11457 => x"80",
         11458 => x"e2",
         11459 => x"05",
         11460 => x"2a",
         11461 => x"59",
         11462 => x"b2",
         11463 => x"9b",
         11464 => x"12",
         11465 => x"2b",
         11466 => x"5e",
         11467 => x"58",
         11468 => x"a4",
         11469 => x"19",
         11470 => x"b8",
         11471 => x"3d",
         11472 => x"b8",
         11473 => x"2e",
         11474 => x"ff",
         11475 => x"0b",
         11476 => x"0c",
         11477 => x"04",
         11478 => x"94",
         11479 => x"98",
         11480 => x"2b",
         11481 => x"98",
         11482 => x"54",
         11483 => x"7e",
         11484 => x"58",
         11485 => x"e4",
         11486 => x"0d",
         11487 => x"3d",
         11488 => x"3d",
         11489 => x"3d",
         11490 => x"80",
         11491 => x"53",
         11492 => x"fd",
         11493 => x"80",
         11494 => x"cf",
         11495 => x"b8",
         11496 => x"84",
         11497 => x"83",
         11498 => x"80",
         11499 => x"7f",
         11500 => x"08",
         11501 => x"0c",
         11502 => x"3d",
         11503 => x"79",
         11504 => x"cc",
         11505 => x"3d",
         11506 => x"5b",
         11507 => x"51",
         11508 => x"3f",
         11509 => x"08",
         11510 => x"e4",
         11511 => x"38",
         11512 => x"3d",
         11513 => x"b4",
         11514 => x"2e",
         11515 => x"b8",
         11516 => x"17",
         11517 => x"7d",
         11518 => x"81",
         11519 => x"b8",
         11520 => x"16",
         11521 => x"8b",
         11522 => x"b8",
         11523 => x"2e",
         11524 => x"57",
         11525 => x"b4",
         11526 => x"82",
         11527 => x"df",
         11528 => x"11",
         11529 => x"33",
         11530 => x"07",
         11531 => x"5d",
         11532 => x"56",
         11533 => x"82",
         11534 => x"80",
         11535 => x"80",
         11536 => x"ff",
         11537 => x"84",
         11538 => x"59",
         11539 => x"08",
         11540 => x"80",
         11541 => x"ff",
         11542 => x"84",
         11543 => x"59",
         11544 => x"08",
         11545 => x"df",
         11546 => x"11",
         11547 => x"33",
         11548 => x"07",
         11549 => x"42",
         11550 => x"56",
         11551 => x"81",
         11552 => x"7a",
         11553 => x"84",
         11554 => x"52",
         11555 => x"a4",
         11556 => x"b8",
         11557 => x"84",
         11558 => x"80",
         11559 => x"38",
         11560 => x"83",
         11561 => x"81",
         11562 => x"e4",
         11563 => x"05",
         11564 => x"ff",
         11565 => x"78",
         11566 => x"33",
         11567 => x"80",
         11568 => x"82",
         11569 => x"17",
         11570 => x"33",
         11571 => x"7c",
         11572 => x"17",
         11573 => x"26",
         11574 => x"76",
         11575 => x"38",
         11576 => x"05",
         11577 => x"80",
         11578 => x"11",
         11579 => x"19",
         11580 => x"58",
         11581 => x"34",
         11582 => x"ff",
         11583 => x"3d",
         11584 => x"58",
         11585 => x"80",
         11586 => x"5a",
         11587 => x"38",
         11588 => x"82",
         11589 => x"0b",
         11590 => x"33",
         11591 => x"83",
         11592 => x"70",
         11593 => x"43",
         11594 => x"5a",
         11595 => x"8d",
         11596 => x"70",
         11597 => x"57",
         11598 => x"f5",
         11599 => x"5b",
         11600 => x"ab",
         11601 => x"76",
         11602 => x"38",
         11603 => x"7e",
         11604 => x"81",
         11605 => x"81",
         11606 => x"77",
         11607 => x"ba",
         11608 => x"05",
         11609 => x"ff",
         11610 => x"06",
         11611 => x"91",
         11612 => x"34",
         11613 => x"e4",
         11614 => x"3d",
         11615 => x"16",
         11616 => x"33",
         11617 => x"71",
         11618 => x"79",
         11619 => x"5e",
         11620 => x"95",
         11621 => x"17",
         11622 => x"2b",
         11623 => x"07",
         11624 => x"dd",
         11625 => x"5d",
         11626 => x"51",
         11627 => x"3f",
         11628 => x"08",
         11629 => x"e4",
         11630 => x"fd",
         11631 => x"b1",
         11632 => x"b4",
         11633 => x"b8",
         11634 => x"81",
         11635 => x"5e",
         11636 => x"3f",
         11637 => x"b8",
         11638 => x"be",
         11639 => x"e4",
         11640 => x"34",
         11641 => x"a8",
         11642 => x"84",
         11643 => x"5a",
         11644 => x"17",
         11645 => x"83",
         11646 => x"33",
         11647 => x"2e",
         11648 => x"fb",
         11649 => x"54",
         11650 => x"a0",
         11651 => x"53",
         11652 => x"16",
         11653 => x"88",
         11654 => x"59",
         11655 => x"ff",
         11656 => x"3d",
         11657 => x"58",
         11658 => x"80",
         11659 => x"c0",
         11660 => x"10",
         11661 => x"05",
         11662 => x"33",
         11663 => x"5e",
         11664 => x"2e",
         11665 => x"fd",
         11666 => x"f1",
         11667 => x"3d",
         11668 => x"19",
         11669 => x"33",
         11670 => x"05",
         11671 => x"60",
         11672 => x"38",
         11673 => x"08",
         11674 => x"59",
         11675 => x"7c",
         11676 => x"5e",
         11677 => x"26",
         11678 => x"f5",
         11679 => x"80",
         11680 => x"84",
         11681 => x"80",
         11682 => x"04",
         11683 => x"7b",
         11684 => x"89",
         11685 => x"2e",
         11686 => x"08",
         11687 => x"2e",
         11688 => x"33",
         11689 => x"2e",
         11690 => x"14",
         11691 => x"22",
         11692 => x"78",
         11693 => x"38",
         11694 => x"5a",
         11695 => x"81",
         11696 => x"15",
         11697 => x"81",
         11698 => x"15",
         11699 => x"76",
         11700 => x"38",
         11701 => x"54",
         11702 => x"78",
         11703 => x"38",
         11704 => x"22",
         11705 => x"52",
         11706 => x"78",
         11707 => x"38",
         11708 => x"17",
         11709 => x"ad",
         11710 => x"e4",
         11711 => x"77",
         11712 => x"55",
         11713 => x"9d",
         11714 => x"e4",
         11715 => x"81",
         11716 => x"30",
         11717 => x"94",
         11718 => x"71",
         11719 => x"08",
         11720 => x"73",
         11721 => x"98",
         11722 => x"27",
         11723 => x"76",
         11724 => x"16",
         11725 => x"17",
         11726 => x"33",
         11727 => x"81",
         11728 => x"57",
         11729 => x"81",
         11730 => x"52",
         11731 => x"99",
         11732 => x"b8",
         11733 => x"84",
         11734 => x"80",
         11735 => x"38",
         11736 => x"98",
         11737 => x"27",
         11738 => x"79",
         11739 => x"14",
         11740 => x"aa",
         11741 => x"16",
         11742 => x"39",
         11743 => x"16",
         11744 => x"72",
         11745 => x"0c",
         11746 => x"04",
         11747 => x"70",
         11748 => x"06",
         11749 => x"fe",
         11750 => x"94",
         11751 => x"57",
         11752 => x"78",
         11753 => x"06",
         11754 => x"77",
         11755 => x"94",
         11756 => x"75",
         11757 => x"38",
         11758 => x"0c",
         11759 => x"80",
         11760 => x"76",
         11761 => x"73",
         11762 => x"59",
         11763 => x"8c",
         11764 => x"08",
         11765 => x"38",
         11766 => x"0c",
         11767 => x"b8",
         11768 => x"3d",
         11769 => x"0b",
         11770 => x"88",
         11771 => x"73",
         11772 => x"fe",
         11773 => x"16",
         11774 => x"2e",
         11775 => x"fe",
         11776 => x"b8",
         11777 => x"94",
         11778 => x"94",
         11779 => x"83",
         11780 => x"75",
         11781 => x"38",
         11782 => x"9c",
         11783 => x"05",
         11784 => x"73",
         11785 => x"f6",
         11786 => x"22",
         11787 => x"b0",
         11788 => x"78",
         11789 => x"5a",
         11790 => x"80",
         11791 => x"38",
         11792 => x"56",
         11793 => x"73",
         11794 => x"ff",
         11795 => x"84",
         11796 => x"54",
         11797 => x"81",
         11798 => x"ff",
         11799 => x"84",
         11800 => x"81",
         11801 => x"fc",
         11802 => x"75",
         11803 => x"fc",
         11804 => x"52",
         11805 => x"97",
         11806 => x"b8",
         11807 => x"84",
         11808 => x"81",
         11809 => x"84",
         11810 => x"ff",
         11811 => x"38",
         11812 => x"08",
         11813 => x"73",
         11814 => x"fe",
         11815 => x"0b",
         11816 => x"82",
         11817 => x"e4",
         11818 => x"0d",
         11819 => x"0d",
         11820 => x"54",
         11821 => x"a2",
         11822 => x"8c",
         11823 => x"52",
         11824 => x"05",
         11825 => x"3f",
         11826 => x"08",
         11827 => x"e4",
         11828 => x"8f",
         11829 => x"0c",
         11830 => x"84",
         11831 => x"8c",
         11832 => x"7a",
         11833 => x"52",
         11834 => x"b9",
         11835 => x"b8",
         11836 => x"84",
         11837 => x"80",
         11838 => x"16",
         11839 => x"2b",
         11840 => x"78",
         11841 => x"86",
         11842 => x"84",
         11843 => x"5b",
         11844 => x"2e",
         11845 => x"9c",
         11846 => x"11",
         11847 => x"33",
         11848 => x"07",
         11849 => x"5d",
         11850 => x"57",
         11851 => x"b3",
         11852 => x"17",
         11853 => x"86",
         11854 => x"17",
         11855 => x"75",
         11856 => x"b9",
         11857 => x"e4",
         11858 => x"84",
         11859 => x"74",
         11860 => x"84",
         11861 => x"0c",
         11862 => x"85",
         11863 => x"0c",
         11864 => x"95",
         11865 => x"18",
         11866 => x"2b",
         11867 => x"07",
         11868 => x"19",
         11869 => x"ff",
         11870 => x"3d",
         11871 => x"89",
         11872 => x"2e",
         11873 => x"08",
         11874 => x"2e",
         11875 => x"33",
         11876 => x"2e",
         11877 => x"13",
         11878 => x"22",
         11879 => x"76",
         11880 => x"80",
         11881 => x"73",
         11882 => x"75",
         11883 => x"b8",
         11884 => x"3d",
         11885 => x"13",
         11886 => x"ff",
         11887 => x"b8",
         11888 => x"06",
         11889 => x"38",
         11890 => x"53",
         11891 => x"f8",
         11892 => x"7c",
         11893 => x"56",
         11894 => x"9f",
         11895 => x"54",
         11896 => x"97",
         11897 => x"53",
         11898 => x"8f",
         11899 => x"22",
         11900 => x"59",
         11901 => x"2e",
         11902 => x"80",
         11903 => x"75",
         11904 => x"c7",
         11905 => x"2e",
         11906 => x"75",
         11907 => x"ff",
         11908 => x"84",
         11909 => x"53",
         11910 => x"08",
         11911 => x"38",
         11912 => x"08",
         11913 => x"52",
         11914 => x"b2",
         11915 => x"52",
         11916 => x"99",
         11917 => x"b8",
         11918 => x"32",
         11919 => x"72",
         11920 => x"84",
         11921 => x"06",
         11922 => x"72",
         11923 => x"0c",
         11924 => x"04",
         11925 => x"75",
         11926 => x"b1",
         11927 => x"52",
         11928 => x"99",
         11929 => x"b8",
         11930 => x"32",
         11931 => x"72",
         11932 => x"84",
         11933 => x"06",
         11934 => x"cf",
         11935 => x"74",
         11936 => x"f9",
         11937 => x"e4",
         11938 => x"e4",
         11939 => x"0d",
         11940 => x"33",
         11941 => x"e8",
         11942 => x"e4",
         11943 => x"53",
         11944 => x"38",
         11945 => x"54",
         11946 => x"39",
         11947 => x"66",
         11948 => x"89",
         11949 => x"97",
         11950 => x"c1",
         11951 => x"b8",
         11952 => x"84",
         11953 => x"80",
         11954 => x"74",
         11955 => x"0c",
         11956 => x"04",
         11957 => x"51",
         11958 => x"3f",
         11959 => x"08",
         11960 => x"e4",
         11961 => x"02",
         11962 => x"33",
         11963 => x"55",
         11964 => x"24",
         11965 => x"80",
         11966 => x"76",
         11967 => x"ff",
         11968 => x"74",
         11969 => x"0c",
         11970 => x"04",
         11971 => x"b8",
         11972 => x"3d",
         11973 => x"3d",
         11974 => x"56",
         11975 => x"95",
         11976 => x"52",
         11977 => x"c0",
         11978 => x"b8",
         11979 => x"84",
         11980 => x"9a",
         11981 => x"0c",
         11982 => x"11",
         11983 => x"94",
         11984 => x"57",
         11985 => x"75",
         11986 => x"75",
         11987 => x"84",
         11988 => x"95",
         11989 => x"84",
         11990 => x"77",
         11991 => x"78",
         11992 => x"93",
         11993 => x"18",
         11994 => x"e4",
         11995 => x"59",
         11996 => x"38",
         11997 => x"71",
         11998 => x"b4",
         11999 => x"2e",
         12000 => x"83",
         12001 => x"5f",
         12002 => x"8d",
         12003 => x"75",
         12004 => x"52",
         12005 => x"51",
         12006 => x"3f",
         12007 => x"08",
         12008 => x"38",
         12009 => x"5e",
         12010 => x"0c",
         12011 => x"57",
         12012 => x"38",
         12013 => x"7d",
         12014 => x"8d",
         12015 => x"b8",
         12016 => x"33",
         12017 => x"71",
         12018 => x"88",
         12019 => x"14",
         12020 => x"07",
         12021 => x"33",
         12022 => x"ff",
         12023 => x"07",
         12024 => x"80",
         12025 => x"60",
         12026 => x"ff",
         12027 => x"05",
         12028 => x"53",
         12029 => x"58",
         12030 => x"78",
         12031 => x"7a",
         12032 => x"94",
         12033 => x"17",
         12034 => x"58",
         12035 => x"34",
         12036 => x"e4",
         12037 => x"0d",
         12038 => x"b4",
         12039 => x"b8",
         12040 => x"81",
         12041 => x"5d",
         12042 => x"3f",
         12043 => x"b8",
         12044 => x"f8",
         12045 => x"e4",
         12046 => x"34",
         12047 => x"a8",
         12048 => x"84",
         12049 => x"5f",
         12050 => x"18",
         12051 => x"bd",
         12052 => x"33",
         12053 => x"2e",
         12054 => x"fe",
         12055 => x"54",
         12056 => x"a0",
         12057 => x"53",
         12058 => x"17",
         12059 => x"fb",
         12060 => x"5e",
         12061 => x"82",
         12062 => x"3d",
         12063 => x"52",
         12064 => x"81",
         12065 => x"b8",
         12066 => x"2e",
         12067 => x"84",
         12068 => x"81",
         12069 => x"38",
         12070 => x"08",
         12071 => x"b8",
         12072 => x"80",
         12073 => x"81",
         12074 => x"58",
         12075 => x"17",
         12076 => x"ca",
         12077 => x"0c",
         12078 => x"0c",
         12079 => x"81",
         12080 => x"84",
         12081 => x"c8",
         12082 => x"b8",
         12083 => x"33",
         12084 => x"88",
         12085 => x"30",
         12086 => x"1f",
         12087 => x"ff",
         12088 => x"5f",
         12089 => x"5f",
         12090 => x"fd",
         12091 => x"8f",
         12092 => x"fd",
         12093 => x"60",
         12094 => x"7f",
         12095 => x"18",
         12096 => x"33",
         12097 => x"77",
         12098 => x"fe",
         12099 => x"60",
         12100 => x"39",
         12101 => x"7b",
         12102 => x"76",
         12103 => x"38",
         12104 => x"74",
         12105 => x"38",
         12106 => x"73",
         12107 => x"38",
         12108 => x"84",
         12109 => x"59",
         12110 => x"81",
         12111 => x"54",
         12112 => x"80",
         12113 => x"17",
         12114 => x"80",
         12115 => x"17",
         12116 => x"2a",
         12117 => x"58",
         12118 => x"80",
         12119 => x"38",
         12120 => x"54",
         12121 => x"08",
         12122 => x"73",
         12123 => x"88",
         12124 => x"08",
         12125 => x"74",
         12126 => x"9c",
         12127 => x"26",
         12128 => x"56",
         12129 => x"18",
         12130 => x"08",
         12131 => x"77",
         12132 => x"59",
         12133 => x"34",
         12134 => x"85",
         12135 => x"18",
         12136 => x"74",
         12137 => x"0c",
         12138 => x"04",
         12139 => x"78",
         12140 => x"38",
         12141 => x"51",
         12142 => x"3f",
         12143 => x"08",
         12144 => x"e4",
         12145 => x"80",
         12146 => x"b8",
         12147 => x"2e",
         12148 => x"84",
         12149 => x"ff",
         12150 => x"38",
         12151 => x"52",
         12152 => x"85",
         12153 => x"b8",
         12154 => x"c8",
         12155 => x"08",
         12156 => x"18",
         12157 => x"58",
         12158 => x"ff",
         12159 => x"15",
         12160 => x"84",
         12161 => x"07",
         12162 => x"17",
         12163 => x"77",
         12164 => x"a0",
         12165 => x"81",
         12166 => x"fe",
         12167 => x"84",
         12168 => x"81",
         12169 => x"fe",
         12170 => x"77",
         12171 => x"fe",
         12172 => x"0b",
         12173 => x"59",
         12174 => x"80",
         12175 => x"0c",
         12176 => x"98",
         12177 => x"76",
         12178 => x"b9",
         12179 => x"e4",
         12180 => x"81",
         12181 => x"b8",
         12182 => x"2e",
         12183 => x"75",
         12184 => x"79",
         12185 => x"e4",
         12186 => x"08",
         12187 => x"38",
         12188 => x"08",
         12189 => x"78",
         12190 => x"54",
         12191 => x"b8",
         12192 => x"81",
         12193 => x"b8",
         12194 => x"17",
         12195 => x"96",
         12196 => x"2e",
         12197 => x"53",
         12198 => x"51",
         12199 => x"3f",
         12200 => x"08",
         12201 => x"e4",
         12202 => x"38",
         12203 => x"51",
         12204 => x"3f",
         12205 => x"08",
         12206 => x"e4",
         12207 => x"80",
         12208 => x"b8",
         12209 => x"2e",
         12210 => x"84",
         12211 => x"ff",
         12212 => x"38",
         12213 => x"52",
         12214 => x"83",
         12215 => x"b8",
         12216 => x"e6",
         12217 => x"08",
         12218 => x"18",
         12219 => x"58",
         12220 => x"90",
         12221 => x"94",
         12222 => x"16",
         12223 => x"54",
         12224 => x"34",
         12225 => x"79",
         12226 => x"38",
         12227 => x"56",
         12228 => x"58",
         12229 => x"81",
         12230 => x"39",
         12231 => x"18",
         12232 => x"fc",
         12233 => x"56",
         12234 => x"0b",
         12235 => x"59",
         12236 => x"39",
         12237 => x"08",
         12238 => x"59",
         12239 => x"39",
         12240 => x"18",
         12241 => x"fd",
         12242 => x"b8",
         12243 => x"c0",
         12244 => x"ff",
         12245 => x"3d",
         12246 => x"a7",
         12247 => x"05",
         12248 => x"51",
         12249 => x"3f",
         12250 => x"08",
         12251 => x"e4",
         12252 => x"8a",
         12253 => x"b8",
         12254 => x"3d",
         12255 => x"4b",
         12256 => x"52",
         12257 => x"52",
         12258 => x"f8",
         12259 => x"e4",
         12260 => x"b8",
         12261 => x"38",
         12262 => x"05",
         12263 => x"2a",
         12264 => x"57",
         12265 => x"cd",
         12266 => x"2b",
         12267 => x"24",
         12268 => x"80",
         12269 => x"70",
         12270 => x"57",
         12271 => x"ff",
         12272 => x"a3",
         12273 => x"11",
         12274 => x"33",
         12275 => x"07",
         12276 => x"5e",
         12277 => x"7c",
         12278 => x"d5",
         12279 => x"2a",
         12280 => x"76",
         12281 => x"ed",
         12282 => x"98",
         12283 => x"2e",
         12284 => x"77",
         12285 => x"84",
         12286 => x"52",
         12287 => x"52",
         12288 => x"f9",
         12289 => x"e4",
         12290 => x"b8",
         12291 => x"e5",
         12292 => x"e4",
         12293 => x"51",
         12294 => x"3f",
         12295 => x"08",
         12296 => x"e4",
         12297 => x"87",
         12298 => x"e4",
         12299 => x"0d",
         12300 => x"33",
         12301 => x"71",
         12302 => x"90",
         12303 => x"07",
         12304 => x"ff",
         12305 => x"b8",
         12306 => x"2e",
         12307 => x"b8",
         12308 => x"a1",
         12309 => x"6f",
         12310 => x"57",
         12311 => x"ff",
         12312 => x"38",
         12313 => x"51",
         12314 => x"3f",
         12315 => x"08",
         12316 => x"e4",
         12317 => x"be",
         12318 => x"70",
         12319 => x"25",
         12320 => x"80",
         12321 => x"74",
         12322 => x"38",
         12323 => x"58",
         12324 => x"27",
         12325 => x"17",
         12326 => x"81",
         12327 => x"56",
         12328 => x"38",
         12329 => x"f5",
         12330 => x"b8",
         12331 => x"b8",
         12332 => x"3d",
         12333 => x"17",
         12334 => x"08",
         12335 => x"b4",
         12336 => x"2e",
         12337 => x"83",
         12338 => x"59",
         12339 => x"2e",
         12340 => x"80",
         12341 => x"54",
         12342 => x"17",
         12343 => x"33",
         12344 => x"ee",
         12345 => x"e4",
         12346 => x"85",
         12347 => x"81",
         12348 => x"18",
         12349 => x"77",
         12350 => x"19",
         12351 => x"78",
         12352 => x"83",
         12353 => x"19",
         12354 => x"fe",
         12355 => x"52",
         12356 => x"8b",
         12357 => x"b8",
         12358 => x"84",
         12359 => x"80",
         12360 => x"38",
         12361 => x"09",
         12362 => x"cd",
         12363 => x"fe",
         12364 => x"54",
         12365 => x"53",
         12366 => x"17",
         12367 => x"f2",
         12368 => x"58",
         12369 => x"08",
         12370 => x"81",
         12371 => x"38",
         12372 => x"08",
         12373 => x"b4",
         12374 => x"18",
         12375 => x"b8",
         12376 => x"55",
         12377 => x"08",
         12378 => x"38",
         12379 => x"55",
         12380 => x"09",
         12381 => x"de",
         12382 => x"b4",
         12383 => x"18",
         12384 => x"7c",
         12385 => x"33",
         12386 => x"c5",
         12387 => x"fe",
         12388 => x"55",
         12389 => x"80",
         12390 => x"52",
         12391 => x"f6",
         12392 => x"b8",
         12393 => x"84",
         12394 => x"80",
         12395 => x"38",
         12396 => x"08",
         12397 => x"e6",
         12398 => x"e4",
         12399 => x"80",
         12400 => x"53",
         12401 => x"51",
         12402 => x"3f",
         12403 => x"08",
         12404 => x"17",
         12405 => x"94",
         12406 => x"5c",
         12407 => x"27",
         12408 => x"81",
         12409 => x"0c",
         12410 => x"81",
         12411 => x"84",
         12412 => x"55",
         12413 => x"ff",
         12414 => x"56",
         12415 => x"79",
         12416 => x"39",
         12417 => x"08",
         12418 => x"39",
         12419 => x"90",
         12420 => x"0d",
         12421 => x"3d",
         12422 => x"52",
         12423 => x"ff",
         12424 => x"84",
         12425 => x"56",
         12426 => x"08",
         12427 => x"38",
         12428 => x"e4",
         12429 => x"0d",
         12430 => x"6f",
         12431 => x"70",
         12432 => x"a6",
         12433 => x"b8",
         12434 => x"84",
         12435 => x"8b",
         12436 => x"84",
         12437 => x"9f",
         12438 => x"84",
         12439 => x"84",
         12440 => x"06",
         12441 => x"80",
         12442 => x"70",
         12443 => x"06",
         12444 => x"56",
         12445 => x"38",
         12446 => x"52",
         12447 => x"52",
         12448 => x"c0",
         12449 => x"e4",
         12450 => x"5c",
         12451 => x"08",
         12452 => x"56",
         12453 => x"08",
         12454 => x"f9",
         12455 => x"e4",
         12456 => x"81",
         12457 => x"81",
         12458 => x"84",
         12459 => x"83",
         12460 => x"5a",
         12461 => x"e2",
         12462 => x"9c",
         12463 => x"05",
         12464 => x"5b",
         12465 => x"8d",
         12466 => x"22",
         12467 => x"b0",
         12468 => x"5c",
         12469 => x"18",
         12470 => x"59",
         12471 => x"57",
         12472 => x"70",
         12473 => x"34",
         12474 => x"74",
         12475 => x"58",
         12476 => x"55",
         12477 => x"81",
         12478 => x"54",
         12479 => x"78",
         12480 => x"33",
         12481 => x"c9",
         12482 => x"e4",
         12483 => x"38",
         12484 => x"dc",
         12485 => x"ff",
         12486 => x"54",
         12487 => x"53",
         12488 => x"53",
         12489 => x"52",
         12490 => x"a5",
         12491 => x"84",
         12492 => x"be",
         12493 => x"e4",
         12494 => x"34",
         12495 => x"a8",
         12496 => x"55",
         12497 => x"08",
         12498 => x"38",
         12499 => x"5b",
         12500 => x"09",
         12501 => x"e1",
         12502 => x"b4",
         12503 => x"18",
         12504 => x"77",
         12505 => x"33",
         12506 => x"e5",
         12507 => x"39",
         12508 => x"7d",
         12509 => x"81",
         12510 => x"b4",
         12511 => x"18",
         12512 => x"ac",
         12513 => x"7c",
         12514 => x"f9",
         12515 => x"e4",
         12516 => x"b8",
         12517 => x"2e",
         12518 => x"84",
         12519 => x"81",
         12520 => x"38",
         12521 => x"08",
         12522 => x"84",
         12523 => x"74",
         12524 => x"fe",
         12525 => x"84",
         12526 => x"fc",
         12527 => x"17",
         12528 => x"94",
         12529 => x"5c",
         12530 => x"27",
         12531 => x"18",
         12532 => x"84",
         12533 => x"07",
         12534 => x"18",
         12535 => x"78",
         12536 => x"a1",
         12537 => x"b8",
         12538 => x"3d",
         12539 => x"17",
         12540 => x"83",
         12541 => x"57",
         12542 => x"78",
         12543 => x"06",
         12544 => x"8b",
         12545 => x"56",
         12546 => x"70",
         12547 => x"34",
         12548 => x"75",
         12549 => x"57",
         12550 => x"18",
         12551 => x"90",
         12552 => x"19",
         12553 => x"75",
         12554 => x"34",
         12555 => x"1a",
         12556 => x"80",
         12557 => x"80",
         12558 => x"d1",
         12559 => x"7c",
         12560 => x"06",
         12561 => x"80",
         12562 => x"77",
         12563 => x"7a",
         12564 => x"34",
         12565 => x"74",
         12566 => x"cc",
         12567 => x"a0",
         12568 => x"1a",
         12569 => x"58",
         12570 => x"81",
         12571 => x"77",
         12572 => x"59",
         12573 => x"56",
         12574 => x"7d",
         12575 => x"80",
         12576 => x"64",
         12577 => x"ff",
         12578 => x"57",
         12579 => x"f2",
         12580 => x"88",
         12581 => x"80",
         12582 => x"75",
         12583 => x"83",
         12584 => x"38",
         12585 => x"0b",
         12586 => x"79",
         12587 => x"96",
         12588 => x"e4",
         12589 => x"b8",
         12590 => x"b6",
         12591 => x"84",
         12592 => x"96",
         12593 => x"b8",
         12594 => x"17",
         12595 => x"98",
         12596 => x"cc",
         12597 => x"34",
         12598 => x"5d",
         12599 => x"34",
         12600 => x"59",
         12601 => x"34",
         12602 => x"79",
         12603 => x"d9",
         12604 => x"90",
         12605 => x"34",
         12606 => x"0b",
         12607 => x"7d",
         12608 => x"80",
         12609 => x"e4",
         12610 => x"84",
         12611 => x"9f",
         12612 => x"76",
         12613 => x"74",
         12614 => x"34",
         12615 => x"57",
         12616 => x"17",
         12617 => x"39",
         12618 => x"5b",
         12619 => x"17",
         12620 => x"2a",
         12621 => x"cd",
         12622 => x"59",
         12623 => x"d8",
         12624 => x"57",
         12625 => x"a1",
         12626 => x"2a",
         12627 => x"18",
         12628 => x"2a",
         12629 => x"18",
         12630 => x"90",
         12631 => x"34",
         12632 => x"0b",
         12633 => x"7d",
         12634 => x"98",
         12635 => x"e4",
         12636 => x"96",
         12637 => x"0d",
         12638 => x"3d",
         12639 => x"5b",
         12640 => x"2e",
         12641 => x"70",
         12642 => x"33",
         12643 => x"56",
         12644 => x"2e",
         12645 => x"74",
         12646 => x"ba",
         12647 => x"38",
         12648 => x"3d",
         12649 => x"52",
         12650 => x"ff",
         12651 => x"84",
         12652 => x"56",
         12653 => x"08",
         12654 => x"38",
         12655 => x"e4",
         12656 => x"0d",
         12657 => x"3d",
         12658 => x"08",
         12659 => x"70",
         12660 => x"9f",
         12661 => x"b8",
         12662 => x"84",
         12663 => x"dc",
         12664 => x"bb",
         12665 => x"a0",
         12666 => x"56",
         12667 => x"a0",
         12668 => x"ae",
         12669 => x"58",
         12670 => x"81",
         12671 => x"77",
         12672 => x"59",
         12673 => x"55",
         12674 => x"99",
         12675 => x"78",
         12676 => x"55",
         12677 => x"05",
         12678 => x"70",
         12679 => x"34",
         12680 => x"74",
         12681 => x"3d",
         12682 => x"51",
         12683 => x"3f",
         12684 => x"08",
         12685 => x"e4",
         12686 => x"38",
         12687 => x"08",
         12688 => x"38",
         12689 => x"b8",
         12690 => x"3d",
         12691 => x"33",
         12692 => x"81",
         12693 => x"57",
         12694 => x"26",
         12695 => x"17",
         12696 => x"06",
         12697 => x"59",
         12698 => x"80",
         12699 => x"7f",
         12700 => x"d4",
         12701 => x"5d",
         12702 => x"5c",
         12703 => x"05",
         12704 => x"70",
         12705 => x"33",
         12706 => x"5a",
         12707 => x"99",
         12708 => x"e0",
         12709 => x"ff",
         12710 => x"ff",
         12711 => x"77",
         12712 => x"38",
         12713 => x"81",
         12714 => x"55",
         12715 => x"9f",
         12716 => x"75",
         12717 => x"81",
         12718 => x"77",
         12719 => x"78",
         12720 => x"30",
         12721 => x"9f",
         12722 => x"5d",
         12723 => x"80",
         12724 => x"81",
         12725 => x"5e",
         12726 => x"24",
         12727 => x"7c",
         12728 => x"5b",
         12729 => x"7b",
         12730 => x"b4",
         12731 => x"0c",
         12732 => x"3d",
         12733 => x"52",
         12734 => x"ff",
         12735 => x"84",
         12736 => x"56",
         12737 => x"08",
         12738 => x"fd",
         12739 => x"aa",
         12740 => x"09",
         12741 => x"ac",
         12742 => x"ff",
         12743 => x"84",
         12744 => x"56",
         12745 => x"08",
         12746 => x"6f",
         12747 => x"8d",
         12748 => x"05",
         12749 => x"58",
         12750 => x"70",
         12751 => x"33",
         12752 => x"05",
         12753 => x"1a",
         12754 => x"38",
         12755 => x"05",
         12756 => x"34",
         12757 => x"70",
         12758 => x"06",
         12759 => x"89",
         12760 => x"07",
         12761 => x"19",
         12762 => x"81",
         12763 => x"34",
         12764 => x"70",
         12765 => x"06",
         12766 => x"80",
         12767 => x"38",
         12768 => x"6b",
         12769 => x"38",
         12770 => x"33",
         12771 => x"71",
         12772 => x"72",
         12773 => x"5c",
         12774 => x"2e",
         12775 => x"fe",
         12776 => x"08",
         12777 => x"56",
         12778 => x"82",
         12779 => x"17",
         12780 => x"29",
         12781 => x"05",
         12782 => x"80",
         12783 => x"38",
         12784 => x"58",
         12785 => x"76",
         12786 => x"83",
         12787 => x"7e",
         12788 => x"81",
         12789 => x"b8",
         12790 => x"17",
         12791 => x"e3",
         12792 => x"b8",
         12793 => x"2e",
         12794 => x"58",
         12795 => x"b4",
         12796 => x"57",
         12797 => x"18",
         12798 => x"fb",
         12799 => x"15",
         12800 => x"ae",
         12801 => x"06",
         12802 => x"70",
         12803 => x"06",
         12804 => x"80",
         12805 => x"7b",
         12806 => x"77",
         12807 => x"34",
         12808 => x"7a",
         12809 => x"81",
         12810 => x"75",
         12811 => x"7d",
         12812 => x"34",
         12813 => x"56",
         12814 => x"18",
         12815 => x"81",
         12816 => x"34",
         12817 => x"3d",
         12818 => x"08",
         12819 => x"74",
         12820 => x"38",
         12821 => x"51",
         12822 => x"3f",
         12823 => x"08",
         12824 => x"e4",
         12825 => x"38",
         12826 => x"98",
         12827 => x"80",
         12828 => x"08",
         12829 => x"38",
         12830 => x"7a",
         12831 => x"7a",
         12832 => x"06",
         12833 => x"81",
         12834 => x"b8",
         12835 => x"16",
         12836 => x"e2",
         12837 => x"b8",
         12838 => x"2e",
         12839 => x"57",
         12840 => x"b4",
         12841 => x"55",
         12842 => x"9c",
         12843 => x"e5",
         12844 => x"0b",
         12845 => x"90",
         12846 => x"27",
         12847 => x"52",
         12848 => x"fc",
         12849 => x"b8",
         12850 => x"84",
         12851 => x"80",
         12852 => x"38",
         12853 => x"84",
         12854 => x"38",
         12855 => x"f9",
         12856 => x"51",
         12857 => x"3f",
         12858 => x"08",
         12859 => x"0c",
         12860 => x"04",
         12861 => x"b8",
         12862 => x"3d",
         12863 => x"18",
         12864 => x"33",
         12865 => x"71",
         12866 => x"78",
         12867 => x"5c",
         12868 => x"84",
         12869 => x"84",
         12870 => x"38",
         12871 => x"08",
         12872 => x"a0",
         12873 => x"b8",
         12874 => x"3d",
         12875 => x"54",
         12876 => x"53",
         12877 => x"16",
         12878 => x"e2",
         12879 => x"58",
         12880 => x"08",
         12881 => x"81",
         12882 => x"38",
         12883 => x"08",
         12884 => x"b4",
         12885 => x"17",
         12886 => x"b8",
         12887 => x"55",
         12888 => x"08",
         12889 => x"38",
         12890 => x"5d",
         12891 => x"09",
         12892 => x"93",
         12893 => x"b4",
         12894 => x"17",
         12895 => x"7b",
         12896 => x"33",
         12897 => x"c9",
         12898 => x"fd",
         12899 => x"54",
         12900 => x"53",
         12901 => x"53",
         12902 => x"52",
         12903 => x"b1",
         12904 => x"84",
         12905 => x"fc",
         12906 => x"b8",
         12907 => x"18",
         12908 => x"08",
         12909 => x"31",
         12910 => x"08",
         12911 => x"a0",
         12912 => x"fc",
         12913 => x"17",
         12914 => x"82",
         12915 => x"06",
         12916 => x"81",
         12917 => x"08",
         12918 => x"05",
         12919 => x"81",
         12920 => x"fe",
         12921 => x"79",
         12922 => x"39",
         12923 => x"02",
         12924 => x"33",
         12925 => x"80",
         12926 => x"56",
         12927 => x"96",
         12928 => x"52",
         12929 => x"ff",
         12930 => x"84",
         12931 => x"56",
         12932 => x"08",
         12933 => x"38",
         12934 => x"e4",
         12935 => x"0d",
         12936 => x"66",
         12937 => x"d0",
         12938 => x"96",
         12939 => x"b8",
         12940 => x"84",
         12941 => x"e0",
         12942 => x"cf",
         12943 => x"a0",
         12944 => x"56",
         12945 => x"74",
         12946 => x"71",
         12947 => x"33",
         12948 => x"74",
         12949 => x"56",
         12950 => x"8b",
         12951 => x"55",
         12952 => x"16",
         12953 => x"fe",
         12954 => x"84",
         12955 => x"84",
         12956 => x"96",
         12957 => x"ec",
         12958 => x"57",
         12959 => x"3d",
         12960 => x"97",
         12961 => x"a1",
         12962 => x"b8",
         12963 => x"84",
         12964 => x"80",
         12965 => x"74",
         12966 => x"0c",
         12967 => x"04",
         12968 => x"52",
         12969 => x"05",
         12970 => x"d8",
         12971 => x"e4",
         12972 => x"b8",
         12973 => x"38",
         12974 => x"05",
         12975 => x"06",
         12976 => x"75",
         12977 => x"84",
         12978 => x"19",
         12979 => x"2b",
         12980 => x"56",
         12981 => x"34",
         12982 => x"55",
         12983 => x"34",
         12984 => x"58",
         12985 => x"34",
         12986 => x"54",
         12987 => x"34",
         12988 => x"0b",
         12989 => x"78",
         12990 => x"88",
         12991 => x"e4",
         12992 => x"e4",
         12993 => x"0d",
         12994 => x"0d",
         12995 => x"5b",
         12996 => x"3d",
         12997 => x"9b",
         12998 => x"a0",
         12999 => x"b8",
         13000 => x"b8",
         13001 => x"70",
         13002 => x"08",
         13003 => x"51",
         13004 => x"80",
         13005 => x"81",
         13006 => x"5a",
         13007 => x"a4",
         13008 => x"70",
         13009 => x"25",
         13010 => x"80",
         13011 => x"38",
         13012 => x"06",
         13013 => x"80",
         13014 => x"38",
         13015 => x"08",
         13016 => x"5a",
         13017 => x"77",
         13018 => x"38",
         13019 => x"7a",
         13020 => x"7a",
         13021 => x"06",
         13022 => x"81",
         13023 => x"b8",
         13024 => x"16",
         13025 => x"dc",
         13026 => x"b8",
         13027 => x"2e",
         13028 => x"57",
         13029 => x"b4",
         13030 => x"57",
         13031 => x"7c",
         13032 => x"58",
         13033 => x"74",
         13034 => x"38",
         13035 => x"74",
         13036 => x"38",
         13037 => x"18",
         13038 => x"11",
         13039 => x"33",
         13040 => x"71",
         13041 => x"81",
         13042 => x"72",
         13043 => x"75",
         13044 => x"62",
         13045 => x"5e",
         13046 => x"76",
         13047 => x"0c",
         13048 => x"04",
         13049 => x"40",
         13050 => x"3d",
         13051 => x"fe",
         13052 => x"84",
         13053 => x"57",
         13054 => x"08",
         13055 => x"8d",
         13056 => x"2e",
         13057 => x"fe",
         13058 => x"7b",
         13059 => x"fe",
         13060 => x"54",
         13061 => x"53",
         13062 => x"53",
         13063 => x"52",
         13064 => x"ad",
         13065 => x"84",
         13066 => x"7a",
         13067 => x"06",
         13068 => x"84",
         13069 => x"83",
         13070 => x"16",
         13071 => x"08",
         13072 => x"e4",
         13073 => x"74",
         13074 => x"27",
         13075 => x"82",
         13076 => x"74",
         13077 => x"81",
         13078 => x"38",
         13079 => x"16",
         13080 => x"08",
         13081 => x"52",
         13082 => x"51",
         13083 => x"3f",
         13084 => x"54",
         13085 => x"16",
         13086 => x"33",
         13087 => x"d2",
         13088 => x"e4",
         13089 => x"fe",
         13090 => x"86",
         13091 => x"74",
         13092 => x"bb",
         13093 => x"e4",
         13094 => x"b8",
         13095 => x"e1",
         13096 => x"e4",
         13097 => x"e4",
         13098 => x"59",
         13099 => x"81",
         13100 => x"57",
         13101 => x"33",
         13102 => x"19",
         13103 => x"27",
         13104 => x"70",
         13105 => x"80",
         13106 => x"80",
         13107 => x"38",
         13108 => x"11",
         13109 => x"57",
         13110 => x"2e",
         13111 => x"e1",
         13112 => x"fd",
         13113 => x"3d",
         13114 => x"a1",
         13115 => x"05",
         13116 => x"51",
         13117 => x"3f",
         13118 => x"08",
         13119 => x"e4",
         13120 => x"38",
         13121 => x"8b",
         13122 => x"a0",
         13123 => x"05",
         13124 => x"15",
         13125 => x"38",
         13126 => x"08",
         13127 => x"81",
         13128 => x"58",
         13129 => x"78",
         13130 => x"38",
         13131 => x"3d",
         13132 => x"81",
         13133 => x"18",
         13134 => x"81",
         13135 => x"7c",
         13136 => x"ff",
         13137 => x"ff",
         13138 => x"a1",
         13139 => x"b5",
         13140 => x"e4",
         13141 => x"dc",
         13142 => x"e4",
         13143 => x"ff",
         13144 => x"80",
         13145 => x"38",
         13146 => x"0b",
         13147 => x"33",
         13148 => x"06",
         13149 => x"78",
         13150 => x"d6",
         13151 => x"78",
         13152 => x"38",
         13153 => x"33",
         13154 => x"06",
         13155 => x"74",
         13156 => x"38",
         13157 => x"09",
         13158 => x"38",
         13159 => x"06",
         13160 => x"a3",
         13161 => x"77",
         13162 => x"38",
         13163 => x"81",
         13164 => x"ff",
         13165 => x"38",
         13166 => x"55",
         13167 => x"81",
         13168 => x"81",
         13169 => x"7b",
         13170 => x"5d",
         13171 => x"a3",
         13172 => x"33",
         13173 => x"06",
         13174 => x"5a",
         13175 => x"fe",
         13176 => x"3d",
         13177 => x"56",
         13178 => x"2e",
         13179 => x"80",
         13180 => x"02",
         13181 => x"79",
         13182 => x"5c",
         13183 => x"2e",
         13184 => x"87",
         13185 => x"5a",
         13186 => x"7d",
         13187 => x"80",
         13188 => x"70",
         13189 => x"ef",
         13190 => x"b8",
         13191 => x"84",
         13192 => x"80",
         13193 => x"74",
         13194 => x"b8",
         13195 => x"3d",
         13196 => x"b5",
         13197 => x"9e",
         13198 => x"b8",
         13199 => x"ff",
         13200 => x"74",
         13201 => x"86",
         13202 => x"b8",
         13203 => x"3d",
         13204 => x"e5",
         13205 => x"fe",
         13206 => x"52",
         13207 => x"f4",
         13208 => x"b8",
         13209 => x"84",
         13210 => x"80",
         13211 => x"80",
         13212 => x"38",
         13213 => x"59",
         13214 => x"70",
         13215 => x"33",
         13216 => x"05",
         13217 => x"15",
         13218 => x"38",
         13219 => x"0b",
         13220 => x"7d",
         13221 => x"ec",
         13222 => x"e4",
         13223 => x"56",
         13224 => x"8a",
         13225 => x"8a",
         13226 => x"ff",
         13227 => x"b8",
         13228 => x"2e",
         13229 => x"fe",
         13230 => x"55",
         13231 => x"fe",
         13232 => x"08",
         13233 => x"52",
         13234 => x"b1",
         13235 => x"e4",
         13236 => x"b8",
         13237 => x"2e",
         13238 => x"81",
         13239 => x"b8",
         13240 => x"19",
         13241 => x"16",
         13242 => x"59",
         13243 => x"77",
         13244 => x"83",
         13245 => x"74",
         13246 => x"81",
         13247 => x"38",
         13248 => x"53",
         13249 => x"81",
         13250 => x"fe",
         13251 => x"84",
         13252 => x"80",
         13253 => x"ff",
         13254 => x"76",
         13255 => x"78",
         13256 => x"38",
         13257 => x"08",
         13258 => x"5a",
         13259 => x"e5",
         13260 => x"38",
         13261 => x"80",
         13262 => x"56",
         13263 => x"2e",
         13264 => x"81",
         13265 => x"81",
         13266 => x"81",
         13267 => x"fe",
         13268 => x"84",
         13269 => x"57",
         13270 => x"08",
         13271 => x"86",
         13272 => x"76",
         13273 => x"bf",
         13274 => x"76",
         13275 => x"a0",
         13276 => x"80",
         13277 => x"05",
         13278 => x"15",
         13279 => x"38",
         13280 => x"0b",
         13281 => x"8b",
         13282 => x"57",
         13283 => x"81",
         13284 => x"76",
         13285 => x"58",
         13286 => x"55",
         13287 => x"fd",
         13288 => x"70",
         13289 => x"33",
         13290 => x"05",
         13291 => x"15",
         13292 => x"38",
         13293 => x"6b",
         13294 => x"34",
         13295 => x"0b",
         13296 => x"7d",
         13297 => x"bc",
         13298 => x"e4",
         13299 => x"ce",
         13300 => x"fe",
         13301 => x"54",
         13302 => x"53",
         13303 => x"18",
         13304 => x"d4",
         13305 => x"b8",
         13306 => x"2e",
         13307 => x"80",
         13308 => x"b8",
         13309 => x"19",
         13310 => x"08",
         13311 => x"31",
         13312 => x"19",
         13313 => x"38",
         13314 => x"55",
         13315 => x"b1",
         13316 => x"e4",
         13317 => x"e8",
         13318 => x"81",
         13319 => x"fe",
         13320 => x"84",
         13321 => x"57",
         13322 => x"08",
         13323 => x"b6",
         13324 => x"39",
         13325 => x"59",
         13326 => x"fd",
         13327 => x"a1",
         13328 => x"b4",
         13329 => x"19",
         13330 => x"7a",
         13331 => x"33",
         13332 => x"fd",
         13333 => x"39",
         13334 => x"60",
         13335 => x"05",
         13336 => x"33",
         13337 => x"89",
         13338 => x"2e",
         13339 => x"08",
         13340 => x"2e",
         13341 => x"33",
         13342 => x"2e",
         13343 => x"15",
         13344 => x"22",
         13345 => x"78",
         13346 => x"38",
         13347 => x"5f",
         13348 => x"38",
         13349 => x"56",
         13350 => x"38",
         13351 => x"81",
         13352 => x"17",
         13353 => x"38",
         13354 => x"70",
         13355 => x"06",
         13356 => x"80",
         13357 => x"38",
         13358 => x"22",
         13359 => x"70",
         13360 => x"57",
         13361 => x"87",
         13362 => x"15",
         13363 => x"30",
         13364 => x"9f",
         13365 => x"e4",
         13366 => x"1c",
         13367 => x"53",
         13368 => x"81",
         13369 => x"38",
         13370 => x"78",
         13371 => x"82",
         13372 => x"56",
         13373 => x"74",
         13374 => x"fe",
         13375 => x"81",
         13376 => x"55",
         13377 => x"75",
         13378 => x"82",
         13379 => x"e4",
         13380 => x"81",
         13381 => x"b8",
         13382 => x"2e",
         13383 => x"84",
         13384 => x"81",
         13385 => x"19",
         13386 => x"2e",
         13387 => x"78",
         13388 => x"06",
         13389 => x"56",
         13390 => x"84",
         13391 => x"90",
         13392 => x"87",
         13393 => x"e4",
         13394 => x"0d",
         13395 => x"33",
         13396 => x"ac",
         13397 => x"e4",
         13398 => x"54",
         13399 => x"38",
         13400 => x"55",
         13401 => x"39",
         13402 => x"81",
         13403 => x"7d",
         13404 => x"80",
         13405 => x"81",
         13406 => x"81",
         13407 => x"38",
         13408 => x"52",
         13409 => x"dd",
         13410 => x"b8",
         13411 => x"84",
         13412 => x"ff",
         13413 => x"81",
         13414 => x"57",
         13415 => x"d7",
         13416 => x"90",
         13417 => x"7b",
         13418 => x"8c",
         13419 => x"18",
         13420 => x"18",
         13421 => x"33",
         13422 => x"5c",
         13423 => x"34",
         13424 => x"fe",
         13425 => x"08",
         13426 => x"7a",
         13427 => x"38",
         13428 => x"94",
         13429 => x"15",
         13430 => x"5d",
         13431 => x"34",
         13432 => x"d6",
         13433 => x"ff",
         13434 => x"5b",
         13435 => x"be",
         13436 => x"fe",
         13437 => x"54",
         13438 => x"ff",
         13439 => x"a1",
         13440 => x"f0",
         13441 => x"0d",
         13442 => x"a5",
         13443 => x"88",
         13444 => x"05",
         13445 => x"5f",
         13446 => x"3d",
         13447 => x"5b",
         13448 => x"2e",
         13449 => x"79",
         13450 => x"5b",
         13451 => x"26",
         13452 => x"ba",
         13453 => x"38",
         13454 => x"75",
         13455 => x"92",
         13456 => x"c0",
         13457 => x"76",
         13458 => x"38",
         13459 => x"84",
         13460 => x"70",
         13461 => x"74",
         13462 => x"38",
         13463 => x"75",
         13464 => x"d8",
         13465 => x"b8",
         13466 => x"40",
         13467 => x"52",
         13468 => x"ce",
         13469 => x"b8",
         13470 => x"ff",
         13471 => x"06",
         13472 => x"57",
         13473 => x"38",
         13474 => x"81",
         13475 => x"57",
         13476 => x"38",
         13477 => x"05",
         13478 => x"79",
         13479 => x"b0",
         13480 => x"e4",
         13481 => x"38",
         13482 => x"80",
         13483 => x"38",
         13484 => x"80",
         13485 => x"38",
         13486 => x"06",
         13487 => x"ff",
         13488 => x"2e",
         13489 => x"80",
         13490 => x"f8",
         13491 => x"80",
         13492 => x"f0",
         13493 => x"7f",
         13494 => x"83",
         13495 => x"89",
         13496 => x"08",
         13497 => x"89",
         13498 => x"4c",
         13499 => x"80",
         13500 => x"38",
         13501 => x"80",
         13502 => x"56",
         13503 => x"74",
         13504 => x"7d",
         13505 => x"df",
         13506 => x"74",
         13507 => x"79",
         13508 => x"be",
         13509 => x"84",
         13510 => x"83",
         13511 => x"83",
         13512 => x"61",
         13513 => x"33",
         13514 => x"07",
         13515 => x"57",
         13516 => x"d5",
         13517 => x"06",
         13518 => x"7d",
         13519 => x"05",
         13520 => x"33",
         13521 => x"80",
         13522 => x"38",
         13523 => x"83",
         13524 => x"12",
         13525 => x"2b",
         13526 => x"07",
         13527 => x"70",
         13528 => x"2b",
         13529 => x"07",
         13530 => x"83",
         13531 => x"12",
         13532 => x"2b",
         13533 => x"07",
         13534 => x"70",
         13535 => x"2b",
         13536 => x"07",
         13537 => x"0c",
         13538 => x"0c",
         13539 => x"44",
         13540 => x"59",
         13541 => x"4b",
         13542 => x"57",
         13543 => x"27",
         13544 => x"93",
         13545 => x"80",
         13546 => x"38",
         13547 => x"70",
         13548 => x"49",
         13549 => x"83",
         13550 => x"87",
         13551 => x"82",
         13552 => x"61",
         13553 => x"66",
         13554 => x"83",
         13555 => x"4a",
         13556 => x"58",
         13557 => x"8a",
         13558 => x"ae",
         13559 => x"2a",
         13560 => x"83",
         13561 => x"56",
         13562 => x"2e",
         13563 => x"77",
         13564 => x"83",
         13565 => x"77",
         13566 => x"70",
         13567 => x"58",
         13568 => x"86",
         13569 => x"27",
         13570 => x"52",
         13571 => x"81",
         13572 => x"b8",
         13573 => x"84",
         13574 => x"b8",
         13575 => x"f5",
         13576 => x"81",
         13577 => x"e4",
         13578 => x"b8",
         13579 => x"71",
         13580 => x"83",
         13581 => x"43",
         13582 => x"89",
         13583 => x"5c",
         13584 => x"1f",
         13585 => x"05",
         13586 => x"05",
         13587 => x"72",
         13588 => x"57",
         13589 => x"2e",
         13590 => x"74",
         13591 => x"90",
         13592 => x"60",
         13593 => x"74",
         13594 => x"f2",
         13595 => x"31",
         13596 => x"53",
         13597 => x"52",
         13598 => x"a9",
         13599 => x"e4",
         13600 => x"83",
         13601 => x"38",
         13602 => x"09",
         13603 => x"dd",
         13604 => x"f5",
         13605 => x"e4",
         13606 => x"ac",
         13607 => x"f9",
         13608 => x"55",
         13609 => x"26",
         13610 => x"74",
         13611 => x"39",
         13612 => x"84",
         13613 => x"9f",
         13614 => x"b8",
         13615 => x"81",
         13616 => x"39",
         13617 => x"b8",
         13618 => x"3d",
         13619 => x"f0",
         13620 => x"33",
         13621 => x"81",
         13622 => x"57",
         13623 => x"26",
         13624 => x"1d",
         13625 => x"06",
         13626 => x"58",
         13627 => x"81",
         13628 => x"0b",
         13629 => x"5f",
         13630 => x"7d",
         13631 => x"70",
         13632 => x"33",
         13633 => x"05",
         13634 => x"9f",
         13635 => x"57",
         13636 => x"89",
         13637 => x"70",
         13638 => x"58",
         13639 => x"18",
         13640 => x"26",
         13641 => x"18",
         13642 => x"06",
         13643 => x"30",
         13644 => x"5a",
         13645 => x"2e",
         13646 => x"85",
         13647 => x"be",
         13648 => x"32",
         13649 => x"72",
         13650 => x"7b",
         13651 => x"4a",
         13652 => x"80",
         13653 => x"1c",
         13654 => x"5c",
         13655 => x"ff",
         13656 => x"56",
         13657 => x"9f",
         13658 => x"53",
         13659 => x"51",
         13660 => x"3f",
         13661 => x"b8",
         13662 => x"b6",
         13663 => x"2a",
         13664 => x"b8",
         13665 => x"56",
         13666 => x"bf",
         13667 => x"8e",
         13668 => x"26",
         13669 => x"74",
         13670 => x"fb",
         13671 => x"56",
         13672 => x"7b",
         13673 => x"ba",
         13674 => x"a3",
         13675 => x"f9",
         13676 => x"81",
         13677 => x"57",
         13678 => x"fd",
         13679 => x"6e",
         13680 => x"46",
         13681 => x"39",
         13682 => x"08",
         13683 => x"9d",
         13684 => x"38",
         13685 => x"81",
         13686 => x"fb",
         13687 => x"57",
         13688 => x"e4",
         13689 => x"0d",
         13690 => x"0c",
         13691 => x"62",
         13692 => x"99",
         13693 => x"60",
         13694 => x"74",
         13695 => x"8e",
         13696 => x"ae",
         13697 => x"61",
         13698 => x"76",
         13699 => x"58",
         13700 => x"55",
         13701 => x"8b",
         13702 => x"a0",
         13703 => x"76",
         13704 => x"58",
         13705 => x"81",
         13706 => x"ff",
         13707 => x"ef",
         13708 => x"05",
         13709 => x"34",
         13710 => x"05",
         13711 => x"8d",
         13712 => x"83",
         13713 => x"4b",
         13714 => x"05",
         13715 => x"2a",
         13716 => x"8f",
         13717 => x"61",
         13718 => x"62",
         13719 => x"30",
         13720 => x"61",
         13721 => x"78",
         13722 => x"06",
         13723 => x"92",
         13724 => x"56",
         13725 => x"ff",
         13726 => x"38",
         13727 => x"ff",
         13728 => x"61",
         13729 => x"74",
         13730 => x"6b",
         13731 => x"34",
         13732 => x"05",
         13733 => x"98",
         13734 => x"61",
         13735 => x"ff",
         13736 => x"34",
         13737 => x"05",
         13738 => x"9c",
         13739 => x"88",
         13740 => x"61",
         13741 => x"7e",
         13742 => x"6b",
         13743 => x"34",
         13744 => x"84",
         13745 => x"84",
         13746 => x"61",
         13747 => x"62",
         13748 => x"f7",
         13749 => x"a7",
         13750 => x"61",
         13751 => x"a1",
         13752 => x"34",
         13753 => x"aa",
         13754 => x"83",
         13755 => x"55",
         13756 => x"05",
         13757 => x"2a",
         13758 => x"97",
         13759 => x"80",
         13760 => x"34",
         13761 => x"05",
         13762 => x"ab",
         13763 => x"ac",
         13764 => x"76",
         13765 => x"58",
         13766 => x"81",
         13767 => x"ff",
         13768 => x"ef",
         13769 => x"fe",
         13770 => x"d5",
         13771 => x"83",
         13772 => x"ff",
         13773 => x"81",
         13774 => x"60",
         13775 => x"fe",
         13776 => x"81",
         13777 => x"e4",
         13778 => x"38",
         13779 => x"62",
         13780 => x"9c",
         13781 => x"57",
         13782 => x"70",
         13783 => x"34",
         13784 => x"74",
         13785 => x"75",
         13786 => x"83",
         13787 => x"38",
         13788 => x"f8",
         13789 => x"2e",
         13790 => x"57",
         13791 => x"76",
         13792 => x"45",
         13793 => x"70",
         13794 => x"34",
         13795 => x"59",
         13796 => x"81",
         13797 => x"76",
         13798 => x"75",
         13799 => x"57",
         13800 => x"66",
         13801 => x"76",
         13802 => x"7a",
         13803 => x"79",
         13804 => x"9d",
         13805 => x"e4",
         13806 => x"38",
         13807 => x"57",
         13808 => x"70",
         13809 => x"34",
         13810 => x"74",
         13811 => x"1b",
         13812 => x"58",
         13813 => x"38",
         13814 => x"40",
         13815 => x"ff",
         13816 => x"56",
         13817 => x"83",
         13818 => x"65",
         13819 => x"26",
         13820 => x"55",
         13821 => x"53",
         13822 => x"51",
         13823 => x"3f",
         13824 => x"08",
         13825 => x"74",
         13826 => x"31",
         13827 => x"db",
         13828 => x"62",
         13829 => x"38",
         13830 => x"83",
         13831 => x"8a",
         13832 => x"62",
         13833 => x"38",
         13834 => x"84",
         13835 => x"83",
         13836 => x"5e",
         13837 => x"38",
         13838 => x"56",
         13839 => x"70",
         13840 => x"34",
         13841 => x"78",
         13842 => x"d5",
         13843 => x"aa",
         13844 => x"83",
         13845 => x"78",
         13846 => x"67",
         13847 => x"81",
         13848 => x"34",
         13849 => x"05",
         13850 => x"84",
         13851 => x"43",
         13852 => x"52",
         13853 => x"fc",
         13854 => x"fe",
         13855 => x"34",
         13856 => x"08",
         13857 => x"07",
         13858 => x"86",
         13859 => x"b8",
         13860 => x"87",
         13861 => x"61",
         13862 => x"34",
         13863 => x"c7",
         13864 => x"61",
         13865 => x"34",
         13866 => x"08",
         13867 => x"05",
         13868 => x"83",
         13869 => x"62",
         13870 => x"64",
         13871 => x"05",
         13872 => x"2a",
         13873 => x"83",
         13874 => x"62",
         13875 => x"7e",
         13876 => x"05",
         13877 => x"78",
         13878 => x"79",
         13879 => x"f1",
         13880 => x"84",
         13881 => x"f7",
         13882 => x"53",
         13883 => x"51",
         13884 => x"3f",
         13885 => x"b8",
         13886 => x"b6",
         13887 => x"e4",
         13888 => x"e4",
         13889 => x"0d",
         13890 => x"0c",
         13891 => x"f9",
         13892 => x"1c",
         13893 => x"5c",
         13894 => x"7a",
         13895 => x"91",
         13896 => x"0b",
         13897 => x"22",
         13898 => x"80",
         13899 => x"74",
         13900 => x"38",
         13901 => x"56",
         13902 => x"17",
         13903 => x"57",
         13904 => x"2e",
         13905 => x"75",
         13906 => x"77",
         13907 => x"fc",
         13908 => x"84",
         13909 => x"10",
         13910 => x"05",
         13911 => x"5e",
         13912 => x"80",
         13913 => x"e4",
         13914 => x"8a",
         13915 => x"fd",
         13916 => x"77",
         13917 => x"38",
         13918 => x"e4",
         13919 => x"e4",
         13920 => x"f5",
         13921 => x"38",
         13922 => x"38",
         13923 => x"5b",
         13924 => x"38",
         13925 => x"c8",
         13926 => x"06",
         13927 => x"2e",
         13928 => x"83",
         13929 => x"39",
         13930 => x"05",
         13931 => x"2a",
         13932 => x"a1",
         13933 => x"90",
         13934 => x"61",
         13935 => x"75",
         13936 => x"76",
         13937 => x"34",
         13938 => x"80",
         13939 => x"05",
         13940 => x"80",
         13941 => x"a1",
         13942 => x"05",
         13943 => x"61",
         13944 => x"34",
         13945 => x"05",
         13946 => x"2a",
         13947 => x"a5",
         13948 => x"90",
         13949 => x"61",
         13950 => x"7c",
         13951 => x"75",
         13952 => x"34",
         13953 => x"05",
         13954 => x"ad",
         13955 => x"61",
         13956 => x"80",
         13957 => x"34",
         13958 => x"05",
         13959 => x"b1",
         13960 => x"61",
         13961 => x"80",
         13962 => x"34",
         13963 => x"80",
         13964 => x"a9",
         13965 => x"05",
         13966 => x"80",
         13967 => x"e4",
         13968 => x"55",
         13969 => x"05",
         13970 => x"70",
         13971 => x"34",
         13972 => x"74",
         13973 => x"cd",
         13974 => x"81",
         13975 => x"76",
         13976 => x"58",
         13977 => x"55",
         13978 => x"f9",
         13979 => x"54",
         13980 => x"52",
         13981 => x"be",
         13982 => x"57",
         13983 => x"08",
         13984 => x"7d",
         13985 => x"05",
         13986 => x"83",
         13987 => x"76",
         13988 => x"e4",
         13989 => x"52",
         13990 => x"bf",
         13991 => x"c3",
         13992 => x"84",
         13993 => x"9f",
         13994 => x"b8",
         13995 => x"f8",
         13996 => x"4a",
         13997 => x"81",
         13998 => x"ff",
         13999 => x"05",
         14000 => x"6a",
         14001 => x"84",
         14002 => x"61",
         14003 => x"ff",
         14004 => x"34",
         14005 => x"05",
         14006 => x"88",
         14007 => x"61",
         14008 => x"ff",
         14009 => x"34",
         14010 => x"7c",
         14011 => x"39",
         14012 => x"1f",
         14013 => x"79",
         14014 => x"d5",
         14015 => x"61",
         14016 => x"75",
         14017 => x"57",
         14018 => x"57",
         14019 => x"60",
         14020 => x"7c",
         14021 => x"5e",
         14022 => x"80",
         14023 => x"81",
         14024 => x"80",
         14025 => x"81",
         14026 => x"80",
         14027 => x"80",
         14028 => x"e4",
         14029 => x"f2",
         14030 => x"05",
         14031 => x"61",
         14032 => x"34",
         14033 => x"83",
         14034 => x"7f",
         14035 => x"7a",
         14036 => x"05",
         14037 => x"2a",
         14038 => x"83",
         14039 => x"7a",
         14040 => x"75",
         14041 => x"05",
         14042 => x"2a",
         14043 => x"83",
         14044 => x"82",
         14045 => x"05",
         14046 => x"83",
         14047 => x"76",
         14048 => x"05",
         14049 => x"83",
         14050 => x"80",
         14051 => x"ff",
         14052 => x"81",
         14053 => x"53",
         14054 => x"51",
         14055 => x"3f",
         14056 => x"1f",
         14057 => x"79",
         14058 => x"a5",
         14059 => x"57",
         14060 => x"39",
         14061 => x"7e",
         14062 => x"80",
         14063 => x"05",
         14064 => x"76",
         14065 => x"38",
         14066 => x"8e",
         14067 => x"54",
         14068 => x"52",
         14069 => x"9a",
         14070 => x"81",
         14071 => x"06",
         14072 => x"3d",
         14073 => x"8d",
         14074 => x"74",
         14075 => x"05",
         14076 => x"17",
         14077 => x"2e",
         14078 => x"77",
         14079 => x"80",
         14080 => x"55",
         14081 => x"76",
         14082 => x"b8",
         14083 => x"3d",
         14084 => x"3d",
         14085 => x"84",
         14086 => x"33",
         14087 => x"8a",
         14088 => x"38",
         14089 => x"56",
         14090 => x"9e",
         14091 => x"08",
         14092 => x"05",
         14093 => x"75",
         14094 => x"55",
         14095 => x"8e",
         14096 => x"18",
         14097 => x"88",
         14098 => x"3d",
         14099 => x"3d",
         14100 => x"74",
         14101 => x"52",
         14102 => x"ff",
         14103 => x"74",
         14104 => x"30",
         14105 => x"9f",
         14106 => x"84",
         14107 => x"1c",
         14108 => x"5a",
         14109 => x"39",
         14110 => x"51",
         14111 => x"ff",
         14112 => x"3d",
         14113 => x"ff",
         14114 => x"3d",
         14115 => x"cc",
         14116 => x"80",
         14117 => x"05",
         14118 => x"15",
         14119 => x"38",
         14120 => x"77",
         14121 => x"2e",
         14122 => x"7c",
         14123 => x"24",
         14124 => x"7d",
         14125 => x"05",
         14126 => x"75",
         14127 => x"55",
         14128 => x"b8",
         14129 => x"18",
         14130 => x"88",
         14131 => x"55",
         14132 => x"9e",
         14133 => x"ff",
         14134 => x"75",
         14135 => x"52",
         14136 => x"ff",
         14137 => x"84",
         14138 => x"86",
         14139 => x"2e",
         14140 => x"0b",
         14141 => x"0c",
         14142 => x"04",
         14143 => x"b0",
         14144 => x"54",
         14145 => x"76",
         14146 => x"9d",
         14147 => x"7b",
         14148 => x"70",
         14149 => x"2a",
         14150 => x"5a",
         14151 => x"a5",
         14152 => x"76",
         14153 => x"3f",
         14154 => x"7d",
         14155 => x"0c",
         14156 => x"04",
         14157 => x"75",
         14158 => x"9a",
         14159 => x"53",
         14160 => x"80",
         14161 => x"38",
         14162 => x"ff",
         14163 => x"84",
         14164 => x"85",
         14165 => x"83",
         14166 => x"27",
         14167 => x"b5",
         14168 => x"06",
         14169 => x"80",
         14170 => x"83",
         14171 => x"51",
         14172 => x"9c",
         14173 => x"70",
         14174 => x"06",
         14175 => x"80",
         14176 => x"38",
         14177 => x"e6",
         14178 => x"22",
         14179 => x"39",
         14180 => x"70",
         14181 => x"84",
         14182 => x"53",
         14183 => x"04",
         14184 => x"02",
         14185 => x"02",
         14186 => x"05",
         14187 => x"80",
         14188 => x"ff",
         14189 => x"70",
         14190 => x"b8",
         14191 => x"3d",
         14192 => x"83",
         14193 => x"81",
         14194 => x"70",
         14195 => x"e9",
         14196 => x"83",
         14197 => x"70",
         14198 => x"e4",
         14199 => x"3d",
         14200 => x"3d",
         14201 => x"70",
         14202 => x"26",
         14203 => x"70",
         14204 => x"06",
         14205 => x"56",
         14206 => x"ff",
         14207 => x"38",
         14208 => x"05",
         14209 => x"71",
         14210 => x"25",
         14211 => x"07",
         14212 => x"53",
         14213 => x"71",
         14214 => x"53",
         14215 => x"88",
         14216 => x"81",
         14217 => x"14",
         14218 => x"76",
         14219 => x"71",
         14220 => x"10",
         14221 => x"82",
         14222 => x"54",
         14223 => x"80",
         14224 => x"26",
         14225 => x"52",
         14226 => x"cb",
         14227 => x"70",
         14228 => x"0c",
         14229 => x"04",
         14230 => x"55",
         14231 => x"71",
         14232 => x"38",
         14233 => x"83",
         14234 => x"54",
         14235 => x"c7",
         14236 => x"83",
         14237 => x"57",
         14238 => x"d3",
         14239 => x"16",
         14240 => x"ff",
         14241 => x"f1",
         14242 => x"70",
         14243 => x"06",
         14244 => x"39",
         14245 => x"83",
         14246 => x"57",
         14247 => x"d0",
         14248 => x"ff",
         14249 => x"51",
         14250 => x"16",
         14251 => x"ff",
         14252 => x"c5",
         14253 => x"70",
         14254 => x"06",
         14255 => x"b9",
         14256 => x"31",
         14257 => x"71",
         14258 => x"ff",
         14259 => x"52",
         14260 => x"39",
         14261 => x"10",
         14262 => x"22",
         14263 => x"ef",
         14264 => x"00",
         14265 => x"ff",
         14266 => x"ff",
         14267 => x"ff",
         14268 => x"00",
         14269 => x"8b",
         14270 => x"80",
         14271 => x"75",
         14272 => x"6a",
         14273 => x"5f",
         14274 => x"54",
         14275 => x"49",
         14276 => x"3e",
         14277 => x"33",
         14278 => x"28",
         14279 => x"1d",
         14280 => x"12",
         14281 => x"07",
         14282 => x"fc",
         14283 => x"f1",
         14284 => x"e6",
         14285 => x"db",
         14286 => x"d0",
         14287 => x"c5",
         14288 => x"ba",
         14289 => x"bf",
         14290 => x"59",
         14291 => x"59",
         14292 => x"59",
         14293 => x"59",
         14294 => x"59",
         14295 => x"59",
         14296 => x"59",
         14297 => x"59",
         14298 => x"59",
         14299 => x"59",
         14300 => x"59",
         14301 => x"59",
         14302 => x"59",
         14303 => x"59",
         14304 => x"59",
         14305 => x"59",
         14306 => x"59",
         14307 => x"59",
         14308 => x"59",
         14309 => x"59",
         14310 => x"59",
         14311 => x"59",
         14312 => x"59",
         14313 => x"59",
         14314 => x"59",
         14315 => x"59",
         14316 => x"59",
         14317 => x"59",
         14318 => x"59",
         14319 => x"59",
         14320 => x"59",
         14321 => x"59",
         14322 => x"59",
         14323 => x"59",
         14324 => x"59",
         14325 => x"59",
         14326 => x"59",
         14327 => x"59",
         14328 => x"59",
         14329 => x"59",
         14330 => x"59",
         14331 => x"59",
         14332 => x"71",
         14333 => x"59",
         14334 => x"59",
         14335 => x"59",
         14336 => x"59",
         14337 => x"59",
         14338 => x"59",
         14339 => x"59",
         14340 => x"59",
         14341 => x"59",
         14342 => x"59",
         14343 => x"59",
         14344 => x"59",
         14345 => x"59",
         14346 => x"59",
         14347 => x"59",
         14348 => x"59",
         14349 => x"07",
         14350 => x"06",
         14351 => x"59",
         14352 => x"8a",
         14353 => x"a8",
         14354 => x"67",
         14355 => x"2c",
         14356 => x"ce",
         14357 => x"59",
         14358 => x"59",
         14359 => x"59",
         14360 => x"59",
         14361 => x"59",
         14362 => x"59",
         14363 => x"59",
         14364 => x"59",
         14365 => x"59",
         14366 => x"59",
         14367 => x"59",
         14368 => x"59",
         14369 => x"59",
         14370 => x"59",
         14371 => x"59",
         14372 => x"59",
         14373 => x"59",
         14374 => x"59",
         14375 => x"59",
         14376 => x"59",
         14377 => x"59",
         14378 => x"59",
         14379 => x"59",
         14380 => x"59",
         14381 => x"59",
         14382 => x"59",
         14383 => x"59",
         14384 => x"59",
         14385 => x"59",
         14386 => x"59",
         14387 => x"59",
         14388 => x"59",
         14389 => x"59",
         14390 => x"59",
         14391 => x"59",
         14392 => x"59",
         14393 => x"59",
         14394 => x"59",
         14395 => x"59",
         14396 => x"59",
         14397 => x"59",
         14398 => x"59",
         14399 => x"59",
         14400 => x"59",
         14401 => x"59",
         14402 => x"59",
         14403 => x"59",
         14404 => x"59",
         14405 => x"59",
         14406 => x"59",
         14407 => x"59",
         14408 => x"59",
         14409 => x"ab",
         14410 => x"70",
         14411 => x"59",
         14412 => x"59",
         14413 => x"59",
         14414 => x"59",
         14415 => x"59",
         14416 => x"59",
         14417 => x"59",
         14418 => x"59",
         14419 => x"63",
         14420 => x"58",
         14421 => x"59",
         14422 => x"41",
         14423 => x"59",
         14424 => x"51",
         14425 => x"47",
         14426 => x"3a",
         14427 => x"12",
         14428 => x"2a",
         14429 => x"36",
         14430 => x"42",
         14431 => x"4e",
         14432 => x"1e",
         14433 => x"86",
         14434 => x"74",
         14435 => x"f0",
         14436 => x"3e",
         14437 => x"10",
         14438 => x"cd",
         14439 => x"8a",
         14440 => x"63",
         14441 => x"ba",
         14442 => x"92",
         14443 => x"01",
         14444 => x"19",
         14445 => x"cd",
         14446 => x"f0",
         14447 => x"fa",
         14448 => x"8a",
         14449 => x"cd",
         14450 => x"cd",
         14451 => x"01",
         14452 => x"92",
         14453 => x"63",
         14454 => x"3e",
         14455 => x"6b",
         14456 => x"84",
         14457 => x"a9",
         14458 => x"ca",
         14459 => x"2b",
         14460 => x"ef",
         14461 => x"44",
         14462 => x"94",
         14463 => x"51",
         14464 => x"51",
         14465 => x"51",
         14466 => x"51",
         14467 => x"51",
         14468 => x"51",
         14469 => x"2a",
         14470 => x"51",
         14471 => x"51",
         14472 => x"51",
         14473 => x"51",
         14474 => x"51",
         14475 => x"51",
         14476 => x"51",
         14477 => x"51",
         14478 => x"51",
         14479 => x"51",
         14480 => x"51",
         14481 => x"51",
         14482 => x"51",
         14483 => x"51",
         14484 => x"51",
         14485 => x"51",
         14486 => x"51",
         14487 => x"51",
         14488 => x"51",
         14489 => x"51",
         14490 => x"51",
         14491 => x"51",
         14492 => x"69",
         14493 => x"57",
         14494 => x"44",
         14495 => x"31",
         14496 => x"5b",
         14497 => x"1f",
         14498 => x"0c",
         14499 => x"74",
         14500 => x"51",
         14501 => x"74",
         14502 => x"fc",
         14503 => x"79",
         14504 => x"a5",
         14505 => x"83",
         14506 => x"ea",
         14507 => x"d8",
         14508 => x"c6",
         14509 => x"b7",
         14510 => x"51",
         14511 => x"5b",
         14512 => x"f7",
         14513 => x"66",
         14514 => x"38",
         14515 => x"8f",
         14516 => x"6c",
         14517 => x"4b",
         14518 => x"21",
         14519 => x"f1",
         14520 => x"78",
         14521 => x"cb",
         14522 => x"ba",
         14523 => x"78",
         14524 => x"78",
         14525 => x"78",
         14526 => x"78",
         14527 => x"78",
         14528 => x"78",
         14529 => x"94",
         14530 => x"a2",
         14531 => x"59",
         14532 => x"78",
         14533 => x"78",
         14534 => x"78",
         14535 => x"78",
         14536 => x"78",
         14537 => x"78",
         14538 => x"78",
         14539 => x"78",
         14540 => x"78",
         14541 => x"78",
         14542 => x"78",
         14543 => x"78",
         14544 => x"78",
         14545 => x"78",
         14546 => x"78",
         14547 => x"78",
         14548 => x"78",
         14549 => x"78",
         14550 => x"78",
         14551 => x"16",
         14552 => x"78",
         14553 => x"78",
         14554 => x"78",
         14555 => x"b9",
         14556 => x"c8",
         14557 => x"6a",
         14558 => x"78",
         14559 => x"78",
         14560 => x"78",
         14561 => x"78",
         14562 => x"4f",
         14563 => x"78",
         14564 => x"32",
         14565 => x"9b",
         14566 => x"10",
         14567 => x"10",
         14568 => x"10",
         14569 => x"10",
         14570 => x"10",
         14571 => x"10",
         14572 => x"eb",
         14573 => x"10",
         14574 => x"10",
         14575 => x"10",
         14576 => x"10",
         14577 => x"10",
         14578 => x"10",
         14579 => x"10",
         14580 => x"10",
         14581 => x"10",
         14582 => x"10",
         14583 => x"10",
         14584 => x"10",
         14585 => x"10",
         14586 => x"10",
         14587 => x"10",
         14588 => x"10",
         14589 => x"10",
         14590 => x"10",
         14591 => x"10",
         14592 => x"10",
         14593 => x"10",
         14594 => x"10",
         14595 => x"ad",
         14596 => x"f5",
         14597 => x"e2",
         14598 => x"cf",
         14599 => x"bd",
         14600 => x"80",
         14601 => x"6d",
         14602 => x"5d",
         14603 => x"10",
         14604 => x"4d",
         14605 => x"3d",
         14606 => x"2b",
         14607 => x"19",
         14608 => x"07",
         14609 => x"78",
         14610 => x"67",
         14611 => x"56",
         14612 => x"3f",
         14613 => x"10",
         14614 => x"89",
         14615 => x"6a",
         14616 => x"c6",
         14617 => x"c6",
         14618 => x"c6",
         14619 => x"c6",
         14620 => x"c6",
         14621 => x"c6",
         14622 => x"c6",
         14623 => x"c6",
         14624 => x"c6",
         14625 => x"c6",
         14626 => x"c6",
         14627 => x"c6",
         14628 => x"c6",
         14629 => x"e8",
         14630 => x"c6",
         14631 => x"c6",
         14632 => x"c6",
         14633 => x"c6",
         14634 => x"c6",
         14635 => x"c6",
         14636 => x"b4",
         14637 => x"c6",
         14638 => x"c6",
         14639 => x"3f",
         14640 => x"c6",
         14641 => x"56",
         14642 => x"c7",
         14643 => x"28",
         14644 => x"d4",
         14645 => x"c1",
         14646 => x"b5",
         14647 => x"aa",
         14648 => x"9f",
         14649 => x"94",
         14650 => x"89",
         14651 => x"7d",
         14652 => x"6f",
         14653 => x"01",
         14654 => x"fd",
         14655 => x"fd",
         14656 => x"49",
         14657 => x"fd",
         14658 => x"fd",
         14659 => x"fd",
         14660 => x"fd",
         14661 => x"fd",
         14662 => x"fd",
         14663 => x"fd",
         14664 => x"fd",
         14665 => x"fd",
         14666 => x"7f",
         14667 => x"0d",
         14668 => x"fd",
         14669 => x"fd",
         14670 => x"fd",
         14671 => x"fd",
         14672 => x"fd",
         14673 => x"fd",
         14674 => x"fd",
         14675 => x"fd",
         14676 => x"fd",
         14677 => x"fd",
         14678 => x"fd",
         14679 => x"fd",
         14680 => x"fd",
         14681 => x"fd",
         14682 => x"fd",
         14683 => x"fd",
         14684 => x"fd",
         14685 => x"fd",
         14686 => x"fd",
         14687 => x"fd",
         14688 => x"fd",
         14689 => x"fd",
         14690 => x"fd",
         14691 => x"fd",
         14692 => x"fd",
         14693 => x"fd",
         14694 => x"fd",
         14695 => x"fd",
         14696 => x"fd",
         14697 => x"fd",
         14698 => x"fd",
         14699 => x"fd",
         14700 => x"fd",
         14701 => x"fd",
         14702 => x"fd",
         14703 => x"fd",
         14704 => x"1d",
         14705 => x"fd",
         14706 => x"fd",
         14707 => x"fd",
         14708 => x"fd",
         14709 => x"17",
         14710 => x"fd",
         14711 => x"fd",
         14712 => x"fd",
         14713 => x"fd",
         14714 => x"fd",
         14715 => x"fd",
         14716 => x"fd",
         14717 => x"fd",
         14718 => x"fd",
         14719 => x"fd",
         14720 => x"2b",
         14721 => x"e1",
         14722 => x"b8",
         14723 => x"b8",
         14724 => x"b8",
         14725 => x"fd",
         14726 => x"e1",
         14727 => x"fd",
         14728 => x"fd",
         14729 => x"ff",
         14730 => x"fd",
         14731 => x"fd",
         14732 => x"16",
         14733 => x"0f",
         14734 => x"fd",
         14735 => x"fd",
         14736 => x"58",
         14737 => x"fd",
         14738 => x"18",
         14739 => x"fd",
         14740 => x"fd",
         14741 => x"17",
         14742 => x"69",
         14743 => x"00",
         14744 => x"63",
         14745 => x"00",
         14746 => x"69",
         14747 => x"00",
         14748 => x"61",
         14749 => x"00",
         14750 => x"65",
         14751 => x"00",
         14752 => x"65",
         14753 => x"00",
         14754 => x"70",
         14755 => x"00",
         14756 => x"66",
         14757 => x"00",
         14758 => x"6d",
         14759 => x"00",
         14760 => x"00",
         14761 => x"00",
         14762 => x"00",
         14763 => x"00",
         14764 => x"00",
         14765 => x"00",
         14766 => x"00",
         14767 => x"6c",
         14768 => x"00",
         14769 => x"00",
         14770 => x"74",
         14771 => x"00",
         14772 => x"65",
         14773 => x"00",
         14774 => x"6f",
         14775 => x"00",
         14776 => x"74",
         14777 => x"00",
         14778 => x"00",
         14779 => x"00",
         14780 => x"73",
         14781 => x"00",
         14782 => x"73",
         14783 => x"00",
         14784 => x"6f",
         14785 => x"00",
         14786 => x"00",
         14787 => x"6e",
         14788 => x"20",
         14789 => x"6f",
         14790 => x"00",
         14791 => x"61",
         14792 => x"65",
         14793 => x"69",
         14794 => x"72",
         14795 => x"74",
         14796 => x"00",
         14797 => x"20",
         14798 => x"79",
         14799 => x"65",
         14800 => x"69",
         14801 => x"2e",
         14802 => x"00",
         14803 => x"75",
         14804 => x"63",
         14805 => x"74",
         14806 => x"6d",
         14807 => x"2e",
         14808 => x"00",
         14809 => x"65",
         14810 => x"20",
         14811 => x"6b",
         14812 => x"00",
         14813 => x"65",
         14814 => x"2c",
         14815 => x"65",
         14816 => x"69",
         14817 => x"63",
         14818 => x"65",
         14819 => x"64",
         14820 => x"00",
         14821 => x"6d",
         14822 => x"61",
         14823 => x"74",
         14824 => x"00",
         14825 => x"63",
         14826 => x"61",
         14827 => x"6c",
         14828 => x"69",
         14829 => x"79",
         14830 => x"6d",
         14831 => x"75",
         14832 => x"6f",
         14833 => x"69",
         14834 => x"00",
         14835 => x"6b",
         14836 => x"74",
         14837 => x"61",
         14838 => x"64",
         14839 => x"00",
         14840 => x"76",
         14841 => x"75",
         14842 => x"72",
         14843 => x"20",
         14844 => x"61",
         14845 => x"2e",
         14846 => x"00",
         14847 => x"69",
         14848 => x"72",
         14849 => x"20",
         14850 => x"74",
         14851 => x"65",
         14852 => x"00",
         14853 => x"65",
         14854 => x"6e",
         14855 => x"20",
         14856 => x"61",
         14857 => x"2e",
         14858 => x"00",
         14859 => x"65",
         14860 => x"72",
         14861 => x"79",
         14862 => x"69",
         14863 => x"2e",
         14864 => x"00",
         14865 => x"65",
         14866 => x"64",
         14867 => x"65",
         14868 => x"00",
         14869 => x"61",
         14870 => x"20",
         14871 => x"65",
         14872 => x"65",
         14873 => x"00",
         14874 => x"70",
         14875 => x"20",
         14876 => x"6e",
         14877 => x"00",
         14878 => x"66",
         14879 => x"20",
         14880 => x"6e",
         14881 => x"00",
         14882 => x"6b",
         14883 => x"74",
         14884 => x"61",
         14885 => x"00",
         14886 => x"65",
         14887 => x"6c",
         14888 => x"72",
         14889 => x"00",
         14890 => x"6b",
         14891 => x"72",
         14892 => x"00",
         14893 => x"63",
         14894 => x"2e",
         14895 => x"00",
         14896 => x"75",
         14897 => x"74",
         14898 => x"25",
         14899 => x"74",
         14900 => x"75",
         14901 => x"74",
         14902 => x"73",
         14903 => x"0a",
         14904 => x"00",
         14905 => x"64",
         14906 => x"00",
         14907 => x"6c",
         14908 => x"00",
         14909 => x"00",
         14910 => x"58",
         14911 => x"00",
         14912 => x"00",
         14913 => x"00",
         14914 => x"00",
         14915 => x"58",
         14916 => x"00",
         14917 => x"20",
         14918 => x"20",
         14919 => x"00",
         14920 => x"00",
         14921 => x"25",
         14922 => x"00",
         14923 => x"30",
         14924 => x"30",
         14925 => x"00",
         14926 => x"32",
         14927 => x"00",
         14928 => x"55",
         14929 => x"65",
         14930 => x"30",
         14931 => x"20",
         14932 => x"25",
         14933 => x"2a",
         14934 => x"00",
         14935 => x"20",
         14936 => x"65",
         14937 => x"70",
         14938 => x"61",
         14939 => x"65",
         14940 => x"00",
         14941 => x"54",
         14942 => x"58",
         14943 => x"74",
         14944 => x"75",
         14945 => x"00",
         14946 => x"54",
         14947 => x"58",
         14948 => x"74",
         14949 => x"75",
         14950 => x"00",
         14951 => x"54",
         14952 => x"58",
         14953 => x"74",
         14954 => x"75",
         14955 => x"00",
         14956 => x"54",
         14957 => x"58",
         14958 => x"74",
         14959 => x"75",
         14960 => x"00",
         14961 => x"54",
         14962 => x"52",
         14963 => x"74",
         14964 => x"75",
         14965 => x"00",
         14966 => x"54",
         14967 => x"44",
         14968 => x"74",
         14969 => x"75",
         14970 => x"00",
         14971 => x"20",
         14972 => x"65",
         14973 => x"70",
         14974 => x"00",
         14975 => x"65",
         14976 => x"6e",
         14977 => x"72",
         14978 => x"00",
         14979 => x"74",
         14980 => x"20",
         14981 => x"74",
         14982 => x"72",
         14983 => x"00",
         14984 => x"62",
         14985 => x"67",
         14986 => x"6d",
         14987 => x"2e",
         14988 => x"00",
         14989 => x"6f",
         14990 => x"63",
         14991 => x"74",
         14992 => x"00",
         14993 => x"5f",
         14994 => x"2e",
         14995 => x"00",
         14996 => x"6c",
         14997 => x"74",
         14998 => x"6e",
         14999 => x"61",
         15000 => x"65",
         15001 => x"20",
         15002 => x"64",
         15003 => x"20",
         15004 => x"61",
         15005 => x"69",
         15006 => x"20",
         15007 => x"75",
         15008 => x"79",
         15009 => x"00",
         15010 => x"00",
         15011 => x"5c",
         15012 => x"00",
         15013 => x"00",
         15014 => x"20",
         15015 => x"6d",
         15016 => x"2e",
         15017 => x"00",
         15018 => x"00",
         15019 => x"00",
         15020 => x"5c",
         15021 => x"25",
         15022 => x"73",
         15023 => x"00",
         15024 => x"64",
         15025 => x"62",
         15026 => x"69",
         15027 => x"2e",
         15028 => x"00",
         15029 => x"74",
         15030 => x"69",
         15031 => x"61",
         15032 => x"69",
         15033 => x"69",
         15034 => x"2e",
         15035 => x"00",
         15036 => x"6c",
         15037 => x"20",
         15038 => x"65",
         15039 => x"25",
         15040 => x"78",
         15041 => x"2e",
         15042 => x"00",
         15043 => x"6c",
         15044 => x"74",
         15045 => x"65",
         15046 => x"6f",
         15047 => x"28",
         15048 => x"2e",
         15049 => x"00",
         15050 => x"63",
         15051 => x"6e",
         15052 => x"6f",
         15053 => x"40",
         15054 => x"38",
         15055 => x"2e",
         15056 => x"00",
         15057 => x"6c",
         15058 => x"30",
         15059 => x"2d",
         15060 => x"00",
         15061 => x"6c",
         15062 => x"30",
         15063 => x"00",
         15064 => x"70",
         15065 => x"6e",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"6c",
         15069 => x"30",
         15070 => x"2d",
         15071 => x"38",
         15072 => x"25",
         15073 => x"29",
         15074 => x"00",
         15075 => x"79",
         15076 => x"2e",
         15077 => x"00",
         15078 => x"6c",
         15079 => x"30",
         15080 => x"00",
         15081 => x"61",
         15082 => x"67",
         15083 => x"2e",
         15084 => x"00",
         15085 => x"70",
         15086 => x"6d",
         15087 => x"00",
         15088 => x"6d",
         15089 => x"74",
         15090 => x"00",
         15091 => x"5c",
         15092 => x"25",
         15093 => x"00",
         15094 => x"6f",
         15095 => x"65",
         15096 => x"75",
         15097 => x"64",
         15098 => x"61",
         15099 => x"74",
         15100 => x"6f",
         15101 => x"73",
         15102 => x"6d",
         15103 => x"64",
         15104 => x"00",
         15105 => x"00",
         15106 => x"25",
         15107 => x"64",
         15108 => x"3a",
         15109 => x"25",
         15110 => x"64",
         15111 => x"00",
         15112 => x"20",
         15113 => x"66",
         15114 => x"72",
         15115 => x"6f",
         15116 => x"00",
         15117 => x"65",
         15118 => x"65",
         15119 => x"6d",
         15120 => x"6d",
         15121 => x"65",
         15122 => x"00",
         15123 => x"72",
         15124 => x"65",
         15125 => x"00",
         15126 => x"20",
         15127 => x"20",
         15128 => x"65",
         15129 => x"65",
         15130 => x"72",
         15131 => x"64",
         15132 => x"73",
         15133 => x"25",
         15134 => x"0a",
         15135 => x"00",
         15136 => x"20",
         15137 => x"20",
         15138 => x"6f",
         15139 => x"53",
         15140 => x"74",
         15141 => x"64",
         15142 => x"73",
         15143 => x"25",
         15144 => x"0a",
         15145 => x"00",
         15146 => x"20",
         15147 => x"63",
         15148 => x"74",
         15149 => x"20",
         15150 => x"72",
         15151 => x"20",
         15152 => x"20",
         15153 => x"25",
         15154 => x"0a",
         15155 => x"00",
         15156 => x"63",
         15157 => x"00",
         15158 => x"20",
         15159 => x"20",
         15160 => x"20",
         15161 => x"20",
         15162 => x"20",
         15163 => x"20",
         15164 => x"20",
         15165 => x"25",
         15166 => x"0a",
         15167 => x"00",
         15168 => x"20",
         15169 => x"74",
         15170 => x"43",
         15171 => x"6b",
         15172 => x"65",
         15173 => x"20",
         15174 => x"20",
         15175 => x"25",
         15176 => x"30",
         15177 => x"48",
         15178 => x"00",
         15179 => x"20",
         15180 => x"68",
         15181 => x"65",
         15182 => x"52",
         15183 => x"43",
         15184 => x"6b",
         15185 => x"65",
         15186 => x"25",
         15187 => x"30",
         15188 => x"48",
         15189 => x"00",
         15190 => x"20",
         15191 => x"41",
         15192 => x"6c",
         15193 => x"20",
         15194 => x"71",
         15195 => x"20",
         15196 => x"20",
         15197 => x"25",
         15198 => x"30",
         15199 => x"48",
         15200 => x"00",
         15201 => x"20",
         15202 => x"00",
         15203 => x"20",
         15204 => x"00",
         15205 => x"20",
         15206 => x"54",
         15207 => x"00",
         15208 => x"20",
         15209 => x"49",
         15210 => x"00",
         15211 => x"20",
         15212 => x"48",
         15213 => x"45",
         15214 => x"53",
         15215 => x"00",
         15216 => x"20",
         15217 => x"52",
         15218 => x"52",
         15219 => x"43",
         15220 => x"6e",
         15221 => x"3d",
         15222 => x"64",
         15223 => x"00",
         15224 => x"20",
         15225 => x"45",
         15226 => x"20",
         15227 => x"54",
         15228 => x"72",
         15229 => x"3d",
         15230 => x"64",
         15231 => x"00",
         15232 => x"20",
         15233 => x"43",
         15234 => x"20",
         15235 => x"44",
         15236 => x"63",
         15237 => x"3d",
         15238 => x"64",
         15239 => x"00",
         15240 => x"20",
         15241 => x"20",
         15242 => x"20",
         15243 => x"25",
         15244 => x"3a",
         15245 => x"58",
         15246 => x"00",
         15247 => x"20",
         15248 => x"4d",
         15249 => x"20",
         15250 => x"25",
         15251 => x"3a",
         15252 => x"58",
         15253 => x"00",
         15254 => x"20",
         15255 => x"4e",
         15256 => x"41",
         15257 => x"25",
         15258 => x"3a",
         15259 => x"58",
         15260 => x"00",
         15261 => x"20",
         15262 => x"41",
         15263 => x"20",
         15264 => x"25",
         15265 => x"3a",
         15266 => x"58",
         15267 => x"00",
         15268 => x"20",
         15269 => x"53",
         15270 => x"4d",
         15271 => x"25",
         15272 => x"3a",
         15273 => x"58",
         15274 => x"00",
         15275 => x"72",
         15276 => x"53",
         15277 => x"63",
         15278 => x"69",
         15279 => x"00",
         15280 => x"6e",
         15281 => x"00",
         15282 => x"6d",
         15283 => x"00",
         15284 => x"6c",
         15285 => x"00",
         15286 => x"69",
         15287 => x"00",
         15288 => x"78",
         15289 => x"00",
         15290 => x"00",
         15291 => x"48",
         15292 => x"00",
         15293 => x"02",
         15294 => x"44",
         15295 => x"00",
         15296 => x"03",
         15297 => x"40",
         15298 => x"00",
         15299 => x"04",
         15300 => x"3c",
         15301 => x"00",
         15302 => x"05",
         15303 => x"38",
         15304 => x"00",
         15305 => x"06",
         15306 => x"34",
         15307 => x"00",
         15308 => x"07",
         15309 => x"30",
         15310 => x"00",
         15311 => x"01",
         15312 => x"2c",
         15313 => x"00",
         15314 => x"08",
         15315 => x"28",
         15316 => x"00",
         15317 => x"0b",
         15318 => x"24",
         15319 => x"00",
         15320 => x"09",
         15321 => x"20",
         15322 => x"00",
         15323 => x"0a",
         15324 => x"1c",
         15325 => x"00",
         15326 => x"0d",
         15327 => x"18",
         15328 => x"00",
         15329 => x"0c",
         15330 => x"14",
         15331 => x"00",
         15332 => x"0e",
         15333 => x"10",
         15334 => x"00",
         15335 => x"0f",
         15336 => x"0c",
         15337 => x"00",
         15338 => x"0f",
         15339 => x"08",
         15340 => x"00",
         15341 => x"10",
         15342 => x"04",
         15343 => x"00",
         15344 => x"11",
         15345 => x"00",
         15346 => x"00",
         15347 => x"12",
         15348 => x"fc",
         15349 => x"00",
         15350 => x"13",
         15351 => x"f8",
         15352 => x"00",
         15353 => x"14",
         15354 => x"f4",
         15355 => x"00",
         15356 => x"15",
         15357 => x"00",
         15358 => x"00",
         15359 => x"00",
         15360 => x"00",
         15361 => x"7e",
         15362 => x"7e",
         15363 => x"7e",
         15364 => x"00",
         15365 => x"7e",
         15366 => x"7e",
         15367 => x"7e",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"6e",
         15380 => x"6f",
         15381 => x"2f",
         15382 => x"61",
         15383 => x"68",
         15384 => x"6f",
         15385 => x"66",
         15386 => x"2c",
         15387 => x"73",
         15388 => x"69",
         15389 => x"00",
         15390 => x"74",
         15391 => x"00",
         15392 => x"74",
         15393 => x"00",
         15394 => x"00",
         15395 => x"6c",
         15396 => x"25",
         15397 => x"00",
         15398 => x"6c",
         15399 => x"74",
         15400 => x"65",
         15401 => x"20",
         15402 => x"20",
         15403 => x"74",
         15404 => x"20",
         15405 => x"65",
         15406 => x"20",
         15407 => x"2e",
         15408 => x"00",
         15409 => x"0a",
         15410 => x"00",
         15411 => x"7e",
         15412 => x"00",
         15413 => x"00",
         15414 => x"00",
         15415 => x"00",
         15416 => x"00",
         15417 => x"30",
         15418 => x"00",
         15419 => x"31",
         15420 => x"00",
         15421 => x"32",
         15422 => x"00",
         15423 => x"33",
         15424 => x"00",
         15425 => x"34",
         15426 => x"00",
         15427 => x"35",
         15428 => x"00",
         15429 => x"37",
         15430 => x"00",
         15431 => x"38",
         15432 => x"00",
         15433 => x"39",
         15434 => x"00",
         15435 => x"30",
         15436 => x"00",
         15437 => x"7e",
         15438 => x"00",
         15439 => x"7e",
         15440 => x"00",
         15441 => x"00",
         15442 => x"7e",
         15443 => x"00",
         15444 => x"7e",
         15445 => x"00",
         15446 => x"64",
         15447 => x"2c",
         15448 => x"25",
         15449 => x"64",
         15450 => x"3a",
         15451 => x"78",
         15452 => x"00",
         15453 => x"64",
         15454 => x"2d",
         15455 => x"25",
         15456 => x"64",
         15457 => x"2c",
         15458 => x"00",
         15459 => x"00",
         15460 => x"64",
         15461 => x"00",
         15462 => x"78",
         15463 => x"00",
         15464 => x"25",
         15465 => x"64",
         15466 => x"00",
         15467 => x"6f",
         15468 => x"43",
         15469 => x"6f",
         15470 => x"00",
         15471 => x"25",
         15472 => x"20",
         15473 => x"78",
         15474 => x"00",
         15475 => x"25",
         15476 => x"20",
         15477 => x"78",
         15478 => x"00",
         15479 => x"25",
         15480 => x"20",
         15481 => x"00",
         15482 => x"74",
         15483 => x"20",
         15484 => x"69",
         15485 => x"2e",
         15486 => x"00",
         15487 => x"00",
         15488 => x"3c",
         15489 => x"7f",
         15490 => x"00",
         15491 => x"3d",
         15492 => x"00",
         15493 => x"00",
         15494 => x"33",
         15495 => x"00",
         15496 => x"4d",
         15497 => x"53",
         15498 => x"00",
         15499 => x"4e",
         15500 => x"20",
         15501 => x"46",
         15502 => x"20",
         15503 => x"00",
         15504 => x"4e",
         15505 => x"20",
         15506 => x"46",
         15507 => x"32",
         15508 => x"00",
         15509 => x"fc",
         15510 => x"00",
         15511 => x"00",
         15512 => x"00",
         15513 => x"07",
         15514 => x"12",
         15515 => x"1c",
         15516 => x"00",
         15517 => x"41",
         15518 => x"80",
         15519 => x"49",
         15520 => x"8f",
         15521 => x"4f",
         15522 => x"55",
         15523 => x"9b",
         15524 => x"9f",
         15525 => x"55",
         15526 => x"a7",
         15527 => x"ab",
         15528 => x"af",
         15529 => x"b3",
         15530 => x"b7",
         15531 => x"bb",
         15532 => x"bf",
         15533 => x"c3",
         15534 => x"c7",
         15535 => x"cb",
         15536 => x"cf",
         15537 => x"d3",
         15538 => x"d7",
         15539 => x"db",
         15540 => x"df",
         15541 => x"e3",
         15542 => x"e7",
         15543 => x"eb",
         15544 => x"ef",
         15545 => x"f3",
         15546 => x"f7",
         15547 => x"fb",
         15548 => x"ff",
         15549 => x"3b",
         15550 => x"2f",
         15551 => x"3a",
         15552 => x"7c",
         15553 => x"00",
         15554 => x"04",
         15555 => x"40",
         15556 => x"00",
         15557 => x"00",
         15558 => x"02",
         15559 => x"08",
         15560 => x"20",
         15561 => x"00",
         15562 => x"fc",
         15563 => x"e2",
         15564 => x"e0",
         15565 => x"e7",
         15566 => x"eb",
         15567 => x"ef",
         15568 => x"ec",
         15569 => x"c5",
         15570 => x"e6",
         15571 => x"f4",
         15572 => x"f2",
         15573 => x"f9",
         15574 => x"d6",
         15575 => x"a2",
         15576 => x"a5",
         15577 => x"92",
         15578 => x"ed",
         15579 => x"fa",
         15580 => x"d1",
         15581 => x"ba",
         15582 => x"10",
         15583 => x"bd",
         15584 => x"a1",
         15585 => x"bb",
         15586 => x"92",
         15587 => x"02",
         15588 => x"61",
         15589 => x"56",
         15590 => x"63",
         15591 => x"57",
         15592 => x"5c",
         15593 => x"10",
         15594 => x"34",
         15595 => x"1c",
         15596 => x"3c",
         15597 => x"5f",
         15598 => x"54",
         15599 => x"66",
         15600 => x"50",
         15601 => x"67",
         15602 => x"64",
         15603 => x"59",
         15604 => x"52",
         15605 => x"6b",
         15606 => x"18",
         15607 => x"88",
         15608 => x"8c",
         15609 => x"80",
         15610 => x"df",
         15611 => x"c0",
         15612 => x"c3",
         15613 => x"c4",
         15614 => x"98",
         15615 => x"b4",
         15616 => x"c6",
         15617 => x"29",
         15618 => x"b1",
         15619 => x"64",
         15620 => x"21",
         15621 => x"48",
         15622 => x"19",
         15623 => x"1a",
         15624 => x"b2",
         15625 => x"a0",
         15626 => x"1a",
         15627 => x"17",
         15628 => x"07",
         15629 => x"01",
         15630 => x"00",
         15631 => x"32",
         15632 => x"39",
         15633 => x"4a",
         15634 => x"79",
         15635 => x"80",
         15636 => x"43",
         15637 => x"82",
         15638 => x"84",
         15639 => x"86",
         15640 => x"87",
         15641 => x"8a",
         15642 => x"8b",
         15643 => x"8e",
         15644 => x"90",
         15645 => x"91",
         15646 => x"94",
         15647 => x"96",
         15648 => x"98",
         15649 => x"3d",
         15650 => x"9c",
         15651 => x"20",
         15652 => x"a0",
         15653 => x"a2",
         15654 => x"a4",
         15655 => x"a6",
         15656 => x"a7",
         15657 => x"aa",
         15658 => x"ac",
         15659 => x"ae",
         15660 => x"af",
         15661 => x"b2",
         15662 => x"b3",
         15663 => x"b5",
         15664 => x"b8",
         15665 => x"ba",
         15666 => x"bc",
         15667 => x"be",
         15668 => x"c0",
         15669 => x"c2",
         15670 => x"c4",
         15671 => x"c4",
         15672 => x"c8",
         15673 => x"ca",
         15674 => x"ca",
         15675 => x"10",
         15676 => x"01",
         15677 => x"de",
         15678 => x"f3",
         15679 => x"f1",
         15680 => x"f4",
         15681 => x"28",
         15682 => x"12",
         15683 => x"09",
         15684 => x"3b",
         15685 => x"3d",
         15686 => x"3f",
         15687 => x"41",
         15688 => x"46",
         15689 => x"53",
         15690 => x"81",
         15691 => x"55",
         15692 => x"8a",
         15693 => x"8f",
         15694 => x"90",
         15695 => x"5d",
         15696 => x"5f",
         15697 => x"61",
         15698 => x"94",
         15699 => x"65",
         15700 => x"67",
         15701 => x"96",
         15702 => x"62",
         15703 => x"6d",
         15704 => x"9c",
         15705 => x"71",
         15706 => x"73",
         15707 => x"9f",
         15708 => x"77",
         15709 => x"79",
         15710 => x"7b",
         15711 => x"64",
         15712 => x"7f",
         15713 => x"81",
         15714 => x"a9",
         15715 => x"85",
         15716 => x"87",
         15717 => x"44",
         15718 => x"b2",
         15719 => x"8d",
         15720 => x"8f",
         15721 => x"91",
         15722 => x"7b",
         15723 => x"fd",
         15724 => x"ff",
         15725 => x"04",
         15726 => x"88",
         15727 => x"8a",
         15728 => x"11",
         15729 => x"02",
         15730 => x"a3",
         15731 => x"08",
         15732 => x"03",
         15733 => x"8e",
         15734 => x"d8",
         15735 => x"f2",
         15736 => x"f9",
         15737 => x"f4",
         15738 => x"f6",
         15739 => x"f7",
         15740 => x"fa",
         15741 => x"30",
         15742 => x"50",
         15743 => x"60",
         15744 => x"8a",
         15745 => x"c1",
         15746 => x"cf",
         15747 => x"c0",
         15748 => x"44",
         15749 => x"26",
         15750 => x"00",
         15751 => x"01",
         15752 => x"00",
         15753 => x"a0",
         15754 => x"00",
         15755 => x"10",
         15756 => x"20",
         15757 => x"30",
         15758 => x"40",
         15759 => x"51",
         15760 => x"59",
         15761 => x"5b",
         15762 => x"5d",
         15763 => x"5f",
         15764 => x"08",
         15765 => x"0e",
         15766 => x"bb",
         15767 => x"c9",
         15768 => x"cb",
         15769 => x"db",
         15770 => x"f9",
         15771 => x"eb",
         15772 => x"fb",
         15773 => x"08",
         15774 => x"08",
         15775 => x"08",
         15776 => x"04",
         15777 => x"b9",
         15778 => x"bc",
         15779 => x"01",
         15780 => x"d0",
         15781 => x"e0",
         15782 => x"e5",
         15783 => x"ec",
         15784 => x"01",
         15785 => x"4e",
         15786 => x"32",
         15787 => x"10",
         15788 => x"01",
         15789 => x"d0",
         15790 => x"30",
         15791 => x"60",
         15792 => x"67",
         15793 => x"75",
         15794 => x"80",
         15795 => x"00",
         15796 => x"41",
         15797 => x"00",
         15798 => x"00",
         15799 => x"58",
         15800 => x"00",
         15801 => x"00",
         15802 => x"00",
         15803 => x"60",
         15804 => x"00",
         15805 => x"00",
         15806 => x"00",
         15807 => x"68",
         15808 => x"00",
         15809 => x"00",
         15810 => x"00",
         15811 => x"70",
         15812 => x"00",
         15813 => x"00",
         15814 => x"00",
         15815 => x"78",
         15816 => x"00",
         15817 => x"00",
         15818 => x"00",
         15819 => x"80",
         15820 => x"00",
         15821 => x"00",
         15822 => x"00",
         15823 => x"88",
         15824 => x"00",
         15825 => x"00",
         15826 => x"00",
         15827 => x"90",
         15828 => x"00",
         15829 => x"00",
         15830 => x"00",
         15831 => x"98",
         15832 => x"00",
         15833 => x"00",
         15834 => x"00",
         15835 => x"a0",
         15836 => x"00",
         15837 => x"00",
         15838 => x"00",
         15839 => x"a4",
         15840 => x"00",
         15841 => x"00",
         15842 => x"00",
         15843 => x"a8",
         15844 => x"00",
         15845 => x"00",
         15846 => x"00",
         15847 => x"ac",
         15848 => x"00",
         15849 => x"00",
         15850 => x"00",
         15851 => x"b0",
         15852 => x"00",
         15853 => x"00",
         15854 => x"00",
         15855 => x"b4",
         15856 => x"00",
         15857 => x"00",
         15858 => x"00",
         15859 => x"b8",
         15860 => x"00",
         15861 => x"00",
         15862 => x"00",
         15863 => x"bc",
         15864 => x"00",
         15865 => x"00",
         15866 => x"00",
         15867 => x"c4",
         15868 => x"00",
         15869 => x"00",
         15870 => x"00",
         15871 => x"c8",
         15872 => x"00",
         15873 => x"00",
         15874 => x"00",
         15875 => x"d0",
         15876 => x"00",
         15877 => x"00",
         15878 => x"00",
         15879 => x"d8",
         15880 => x"00",
         15881 => x"00",
         15882 => x"00",
         15883 => x"e0",
         15884 => x"00",
         15885 => x"00",
         15886 => x"00",
         15887 => x"e8",
         15888 => x"00",
         15889 => x"00",
         15890 => x"00",
         15891 => x"ec",
         15892 => x"00",
         15893 => x"00",
         15894 => x"00",
         15895 => x"f0",
         15896 => x"00",
         15897 => x"00",
         15898 => x"00",
         15899 => x"f8",
         15900 => x"00",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"00",
         15905 => x"00",
         15906 => x"00",
         15907 => x"08",
         15908 => x"00",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"ff",
         15914 => x"00",
         15915 => x"ff",
         15916 => x"00",
         15917 => x"ff",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"ff",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"00",
         15926 => x"00",
         15927 => x"00",
         15928 => x"00",
         15929 => x"00",
         15930 => x"01",
         15931 => x"01",
         15932 => x"01",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"78",
         15959 => x"00",
         15960 => x"80",
         15961 => x"00",
         15962 => x"88",
         15963 => x"00",
         15964 => x"80",
         15965 => x"fd",
         15966 => x"0d",
         15967 => x"5b",
         15968 => x"f0",
         15969 => x"74",
         15970 => x"78",
         15971 => x"6c",
         15972 => x"70",
         15973 => x"64",
         15974 => x"68",
         15975 => x"34",
         15976 => x"38",
         15977 => x"20",
         15978 => x"2e",
         15979 => x"f4",
         15980 => x"2f",
         15981 => x"f0",
         15982 => x"f0",
         15983 => x"83",
         15984 => x"f0",
         15985 => x"fd",
         15986 => x"0d",
         15987 => x"5b",
         15988 => x"f0",
         15989 => x"54",
         15990 => x"58",
         15991 => x"4c",
         15992 => x"50",
         15993 => x"44",
         15994 => x"48",
         15995 => x"34",
         15996 => x"38",
         15997 => x"20",
         15998 => x"2e",
         15999 => x"f4",
         16000 => x"2f",
         16001 => x"f0",
         16002 => x"f0",
         16003 => x"83",
         16004 => x"f0",
         16005 => x"fd",
         16006 => x"0d",
         16007 => x"7b",
         16008 => x"f0",
         16009 => x"54",
         16010 => x"58",
         16011 => x"4c",
         16012 => x"50",
         16013 => x"44",
         16014 => x"48",
         16015 => x"24",
         16016 => x"28",
         16017 => x"20",
         16018 => x"3e",
         16019 => x"e1",
         16020 => x"2f",
         16021 => x"f0",
         16022 => x"f0",
         16023 => x"88",
         16024 => x"f0",
         16025 => x"fa",
         16026 => x"f0",
         16027 => x"1b",
         16028 => x"f0",
         16029 => x"14",
         16030 => x"18",
         16031 => x"0c",
         16032 => x"10",
         16033 => x"04",
         16034 => x"08",
         16035 => x"f0",
         16036 => x"f0",
         16037 => x"f0",
         16038 => x"f0",
         16039 => x"f0",
         16040 => x"1c",
         16041 => x"f0",
         16042 => x"f0",
         16043 => x"83",
         16044 => x"f0",
         16045 => x"c9",
         16046 => x"cd",
         16047 => x"b3",
         16048 => x"f0",
         16049 => x"31",
         16050 => x"dd",
         16051 => x"56",
         16052 => x"b1",
         16053 => x"48",
         16054 => x"73",
         16055 => x"3b",
         16056 => x"a2",
         16057 => x"00",
         16058 => x"b9",
         16059 => x"c1",
         16060 => x"be",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"83",
         16064 => x"f0",
         16065 => x"00",
         16066 => x"00",
         16067 => x"00",
         16068 => x"00",
         16069 => x"00",
         16070 => x"00",
         16071 => x"00",
         16072 => x"00",
         16073 => x"00",
         16074 => x"00",
         16075 => x"00",
         16076 => x"00",
         16077 => x"00",
         16078 => x"00",
         16079 => x"00",
         16080 => x"00",
         16081 => x"00",
         16082 => x"00",
         16083 => x"00",
         16084 => x"00",
         16085 => x"00",
         16086 => x"00",
         16087 => x"00",
         16088 => x"00",
         16089 => x"00",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"cc",
         16094 => x"00",
         16095 => x"d4",
         16096 => x"00",
         16097 => x"d8",
         16098 => x"00",
         16099 => x"dc",
         16100 => x"00",
         16101 => x"e0",
         16102 => x"00",
         16103 => x"e4",
         16104 => x"00",
         16105 => x"ec",
         16106 => x"00",
         16107 => x"f4",
         16108 => x"00",
         16109 => x"fc",
         16110 => x"00",
         16111 => x"04",
         16112 => x"00",
         16113 => x"0c",
         16114 => x"00",
         16115 => x"14",
         16116 => x"00",
         16117 => x"1c",
         16118 => x"00",
         16119 => x"24",
         16120 => x"00",
         16121 => x"2c",
         16122 => x"00",
         16123 => x"34",
         16124 => x"00",
         16125 => x"3c",
         16126 => x"00",
         16127 => x"44",
         16128 => x"00",
         16129 => x"48",
         16130 => x"00",
         16131 => x"50",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"19",
         18134 => x"00",
         18135 => x"00",
         18136 => x"f3",
         18137 => x"f7",
         18138 => x"fb",
         18139 => x"ff",
         18140 => x"c3",
         18141 => x"e2",
         18142 => x"e6",
         18143 => x"f4",
         18144 => x"63",
         18145 => x"67",
         18146 => x"6a",
         18147 => x"2d",
         18148 => x"23",
         18149 => x"27",
         18150 => x"2c",
         18151 => x"49",
         18152 => x"03",
         18153 => x"07",
         18154 => x"0b",
         18155 => x"0f",
         18156 => x"13",
         18157 => x"17",
         18158 => x"52",
         18159 => x"3c",
         18160 => x"83",
         18161 => x"87",
         18162 => x"8b",
         18163 => x"8f",
         18164 => x"93",
         18165 => x"97",
         18166 => x"bc",
         18167 => x"c0",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"03",
         18199 => x"01",
         18200 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"e9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"83",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a6",
           270 => x"0b",
           271 => x"0b",
           272 => x"c6",
           273 => x"0b",
           274 => x"0b",
           275 => x"e6",
           276 => x"0b",
           277 => x"0b",
           278 => x"86",
           279 => x"0b",
           280 => x"0b",
           281 => x"a6",
           282 => x"0b",
           283 => x"0b",
           284 => x"c6",
           285 => x"0b",
           286 => x"0b",
           287 => x"e8",
           288 => x"0b",
           289 => x"0b",
           290 => x"8a",
           291 => x"0b",
           292 => x"0b",
           293 => x"ac",
           294 => x"0b",
           295 => x"0b",
           296 => x"ce",
           297 => x"0b",
           298 => x"0b",
           299 => x"f0",
           300 => x"0b",
           301 => x"0b",
           302 => x"92",
           303 => x"0b",
           304 => x"0b",
           305 => x"b4",
           306 => x"0b",
           307 => x"0b",
           308 => x"d6",
           309 => x"0b",
           310 => x"0b",
           311 => x"f8",
           312 => x"0b",
           313 => x"0b",
           314 => x"9a",
           315 => x"0b",
           316 => x"0b",
           317 => x"bc",
           318 => x"0b",
           319 => x"0b",
           320 => x"de",
           321 => x"0b",
           322 => x"0b",
           323 => x"80",
           324 => x"0b",
           325 => x"0b",
           326 => x"a2",
           327 => x"0b",
           328 => x"0b",
           329 => x"c4",
           330 => x"0b",
           331 => x"0b",
           332 => x"e6",
           333 => x"0b",
           334 => x"0b",
           335 => x"88",
           336 => x"0b",
           337 => x"0b",
           338 => x"aa",
           339 => x"0b",
           340 => x"0b",
           341 => x"cb",
           342 => x"0b",
           343 => x"0b",
           344 => x"ed",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"b8",
           386 => x"d5",
           387 => x"b8",
           388 => x"c0",
           389 => x"84",
           390 => x"a2",
           391 => x"b8",
           392 => x"c0",
           393 => x"84",
           394 => x"a0",
           395 => x"b8",
           396 => x"c0",
           397 => x"84",
           398 => x"a0",
           399 => x"b8",
           400 => x"c0",
           401 => x"84",
           402 => x"94",
           403 => x"b8",
           404 => x"c0",
           405 => x"84",
           406 => x"a1",
           407 => x"b8",
           408 => x"c0",
           409 => x"84",
           410 => x"af",
           411 => x"b8",
           412 => x"c0",
           413 => x"84",
           414 => x"ad",
           415 => x"b8",
           416 => x"c0",
           417 => x"84",
           418 => x"94",
           419 => x"b8",
           420 => x"c0",
           421 => x"84",
           422 => x"95",
           423 => x"b8",
           424 => x"c0",
           425 => x"84",
           426 => x"95",
           427 => x"b8",
           428 => x"c0",
           429 => x"84",
           430 => x"b1",
           431 => x"b8",
           432 => x"c0",
           433 => x"84",
           434 => x"80",
           435 => x"84",
           436 => x"80",
           437 => x"04",
           438 => x"0c",
           439 => x"2d",
           440 => x"08",
           441 => x"90",
           442 => x"f0",
           443 => x"8d",
           444 => x"f0",
           445 => x"80",
           446 => x"b8",
           447 => x"d3",
           448 => x"b8",
           449 => x"c0",
           450 => x"84",
           451 => x"82",
           452 => x"84",
           453 => x"80",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"90",
           459 => x"f0",
           460 => x"8d",
           461 => x"f0",
           462 => x"80",
           463 => x"b8",
           464 => x"d7",
           465 => x"b8",
           466 => x"c0",
           467 => x"84",
           468 => x"82",
           469 => x"84",
           470 => x"80",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"90",
           476 => x"f0",
           477 => x"f6",
           478 => x"f0",
           479 => x"80",
           480 => x"b8",
           481 => x"f1",
           482 => x"b8",
           483 => x"c0",
           484 => x"84",
           485 => x"82",
           486 => x"84",
           487 => x"80",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"90",
           493 => x"f0",
           494 => x"91",
           495 => x"f0",
           496 => x"80",
           497 => x"b8",
           498 => x"fe",
           499 => x"b8",
           500 => x"c0",
           501 => x"84",
           502 => x"83",
           503 => x"84",
           504 => x"80",
           505 => x"04",
           506 => x"0c",
           507 => x"2d",
           508 => x"08",
           509 => x"90",
           510 => x"f0",
           511 => x"ec",
           512 => x"f0",
           513 => x"80",
           514 => x"b8",
           515 => x"94",
           516 => x"b8",
           517 => x"c0",
           518 => x"84",
           519 => x"82",
           520 => x"84",
           521 => x"80",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"90",
           527 => x"f0",
           528 => x"fd",
           529 => x"f0",
           530 => x"80",
           531 => x"b8",
           532 => x"f6",
           533 => x"b8",
           534 => x"c0",
           535 => x"84",
           536 => x"83",
           537 => x"84",
           538 => x"80",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"90",
           544 => x"f0",
           545 => x"d8",
           546 => x"f0",
           547 => x"80",
           548 => x"b8",
           549 => x"c6",
           550 => x"b8",
           551 => x"c0",
           552 => x"84",
           553 => x"83",
           554 => x"84",
           555 => x"80",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"90",
           561 => x"f0",
           562 => x"b4",
           563 => x"f0",
           564 => x"80",
           565 => x"b8",
           566 => x"f3",
           567 => x"b8",
           568 => x"c0",
           569 => x"84",
           570 => x"81",
           571 => x"84",
           572 => x"80",
           573 => x"04",
           574 => x"0c",
           575 => x"2d",
           576 => x"08",
           577 => x"90",
           578 => x"f0",
           579 => x"8f",
           580 => x"f0",
           581 => x"80",
           582 => x"b8",
           583 => x"d1",
           584 => x"b8",
           585 => x"c0",
           586 => x"84",
           587 => x"80",
           588 => x"84",
           589 => x"80",
           590 => x"04",
           591 => x"0c",
           592 => x"84",
           593 => x"80",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"90",
           599 => x"f0",
           600 => x"ab",
           601 => x"f0",
           602 => x"80",
           603 => x"b8",
           604 => x"f1",
           605 => x"b8",
           606 => x"c0",
           607 => x"84",
           608 => x"81",
           609 => x"84",
           610 => x"80",
           611 => x"04",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"04",
           621 => x"81",
           622 => x"83",
           623 => x"05",
           624 => x"10",
           625 => x"72",
           626 => x"51",
           627 => x"72",
           628 => x"06",
           629 => x"72",
           630 => x"10",
           631 => x"10",
           632 => x"ed",
           633 => x"53",
           634 => x"b8",
           635 => x"d4",
           636 => x"38",
           637 => x"84",
           638 => x"0b",
           639 => x"ec",
           640 => x"51",
           641 => x"04",
           642 => x"0d",
           643 => x"70",
           644 => x"08",
           645 => x"52",
           646 => x"08",
           647 => x"3f",
           648 => x"04",
           649 => x"78",
           650 => x"11",
           651 => x"81",
           652 => x"25",
           653 => x"55",
           654 => x"72",
           655 => x"81",
           656 => x"38",
           657 => x"74",
           658 => x"30",
           659 => x"9f",
           660 => x"55",
           661 => x"74",
           662 => x"71",
           663 => x"38",
           664 => x"fa",
           665 => x"e4",
           666 => x"b8",
           667 => x"2e",
           668 => x"b8",
           669 => x"70",
           670 => x"34",
           671 => x"8a",
           672 => x"70",
           673 => x"2a",
           674 => x"54",
           675 => x"cb",
           676 => x"34",
           677 => x"84",
           678 => x"88",
           679 => x"80",
           680 => x"e4",
           681 => x"0d",
           682 => x"0d",
           683 => x"02",
           684 => x"05",
           685 => x"fe",
           686 => x"3d",
           687 => x"7e",
           688 => x"e4",
           689 => x"3f",
           690 => x"80",
           691 => x"3d",
           692 => x"3d",
           693 => x"88",
           694 => x"52",
           695 => x"3f",
           696 => x"04",
           697 => x"61",
           698 => x"5d",
           699 => x"8c",
           700 => x"1e",
           701 => x"2a",
           702 => x"06",
           703 => x"ff",
           704 => x"2e",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"81",
           709 => x"06",
           710 => x"80",
           711 => x"38",
           712 => x"7e",
           713 => x"a3",
           714 => x"32",
           715 => x"80",
           716 => x"55",
           717 => x"72",
           718 => x"38",
           719 => x"70",
           720 => x"06",
           721 => x"80",
           722 => x"7a",
           723 => x"5b",
           724 => x"76",
           725 => x"8c",
           726 => x"73",
           727 => x"0c",
           728 => x"04",
           729 => x"54",
           730 => x"10",
           731 => x"70",
           732 => x"98",
           733 => x"81",
           734 => x"8b",
           735 => x"98",
           736 => x"5b",
           737 => x"79",
           738 => x"38",
           739 => x"53",
           740 => x"38",
           741 => x"58",
           742 => x"f7",
           743 => x"39",
           744 => x"09",
           745 => x"38",
           746 => x"5a",
           747 => x"7c",
           748 => x"76",
           749 => x"ff",
           750 => x"52",
           751 => x"af",
           752 => x"57",
           753 => x"38",
           754 => x"7a",
           755 => x"81",
           756 => x"78",
           757 => x"70",
           758 => x"54",
           759 => x"e0",
           760 => x"80",
           761 => x"38",
           762 => x"83",
           763 => x"54",
           764 => x"73",
           765 => x"59",
           766 => x"27",
           767 => x"52",
           768 => x"eb",
           769 => x"33",
           770 => x"fe",
           771 => x"c7",
           772 => x"59",
           773 => x"88",
           774 => x"84",
           775 => x"7d",
           776 => x"06",
           777 => x"54",
           778 => x"5e",
           779 => x"51",
           780 => x"84",
           781 => x"81",
           782 => x"b8",
           783 => x"df",
           784 => x"72",
           785 => x"38",
           786 => x"08",
           787 => x"74",
           788 => x"05",
           789 => x"52",
           790 => x"ca",
           791 => x"e4",
           792 => x"b8",
           793 => x"38",
           794 => x"f4",
           795 => x"7b",
           796 => x"56",
           797 => x"8f",
           798 => x"80",
           799 => x"80",
           800 => x"90",
           801 => x"7a",
           802 => x"81",
           803 => x"73",
           804 => x"38",
           805 => x"80",
           806 => x"80",
           807 => x"90",
           808 => x"77",
           809 => x"29",
           810 => x"05",
           811 => x"2c",
           812 => x"2a",
           813 => x"54",
           814 => x"2e",
           815 => x"98",
           816 => x"ff",
           817 => x"78",
           818 => x"cc",
           819 => x"ff",
           820 => x"83",
           821 => x"2a",
           822 => x"74",
           823 => x"73",
           824 => x"f0",
           825 => x"31",
           826 => x"90",
           827 => x"80",
           828 => x"53",
           829 => x"85",
           830 => x"81",
           831 => x"54",
           832 => x"38",
           833 => x"81",
           834 => x"86",
           835 => x"85",
           836 => x"54",
           837 => x"38",
           838 => x"54",
           839 => x"38",
           840 => x"81",
           841 => x"80",
           842 => x"77",
           843 => x"80",
           844 => x"80",
           845 => x"2c",
           846 => x"80",
           847 => x"38",
           848 => x"51",
           849 => x"77",
           850 => x"80",
           851 => x"80",
           852 => x"2c",
           853 => x"73",
           854 => x"38",
           855 => x"53",
           856 => x"b2",
           857 => x"81",
           858 => x"81",
           859 => x"70",
           860 => x"55",
           861 => x"25",
           862 => x"52",
           863 => x"ef",
           864 => x"81",
           865 => x"81",
           866 => x"70",
           867 => x"55",
           868 => x"24",
           869 => x"87",
           870 => x"06",
           871 => x"80",
           872 => x"38",
           873 => x"2e",
           874 => x"76",
           875 => x"81",
           876 => x"80",
           877 => x"e2",
           878 => x"b8",
           879 => x"38",
           880 => x"1e",
           881 => x"5e",
           882 => x"7d",
           883 => x"2e",
           884 => x"ec",
           885 => x"06",
           886 => x"2e",
           887 => x"77",
           888 => x"80",
           889 => x"80",
           890 => x"2c",
           891 => x"80",
           892 => x"91",
           893 => x"a0",
           894 => x"3f",
           895 => x"90",
           896 => x"a0",
           897 => x"58",
           898 => x"87",
           899 => x"39",
           900 => x"07",
           901 => x"57",
           902 => x"84",
           903 => x"7e",
           904 => x"06",
           905 => x"55",
           906 => x"39",
           907 => x"05",
           908 => x"0a",
           909 => x"33",
           910 => x"72",
           911 => x"80",
           912 => x"80",
           913 => x"90",
           914 => x"5a",
           915 => x"5f",
           916 => x"70",
           917 => x"55",
           918 => x"38",
           919 => x"80",
           920 => x"80",
           921 => x"90",
           922 => x"5f",
           923 => x"fe",
           924 => x"52",
           925 => x"f7",
           926 => x"ff",
           927 => x"ff",
           928 => x"57",
           929 => x"ff",
           930 => x"38",
           931 => x"70",
           932 => x"33",
           933 => x"3f",
           934 => x"1a",
           935 => x"ff",
           936 => x"79",
           937 => x"2e",
           938 => x"7c",
           939 => x"81",
           940 => x"51",
           941 => x"e2",
           942 => x"0a",
           943 => x"0a",
           944 => x"80",
           945 => x"80",
           946 => x"90",
           947 => x"56",
           948 => x"87",
           949 => x"06",
           950 => x"7a",
           951 => x"fe",
           952 => x"60",
           953 => x"08",
           954 => x"41",
           955 => x"24",
           956 => x"7a",
           957 => x"06",
           958 => x"f4",
           959 => x"39",
           960 => x"7c",
           961 => x"76",
           962 => x"f8",
           963 => x"88",
           964 => x"7c",
           965 => x"76",
           966 => x"f8",
           967 => x"60",
           968 => x"08",
           969 => x"56",
           970 => x"72",
           971 => x"75",
           972 => x"3f",
           973 => x"08",
           974 => x"06",
           975 => x"90",
           976 => x"72",
           977 => x"fe",
           978 => x"80",
           979 => x"33",
           980 => x"f7",
           981 => x"ff",
           982 => x"84",
           983 => x"77",
           984 => x"58",
           985 => x"81",
           986 => x"51",
           987 => x"84",
           988 => x"83",
           989 => x"78",
           990 => x"2b",
           991 => x"39",
           992 => x"07",
           993 => x"5b",
           994 => x"38",
           995 => x"77",
           996 => x"80",
           997 => x"80",
           998 => x"2c",
           999 => x"80",
          1000 => x"d6",
          1001 => x"a0",
          1002 => x"3f",
          1003 => x"52",
          1004 => x"bb",
          1005 => x"2e",
          1006 => x"fa",
          1007 => x"52",
          1008 => x"ab",
          1009 => x"2a",
          1010 => x"7e",
          1011 => x"8c",
          1012 => x"39",
          1013 => x"78",
          1014 => x"2b",
          1015 => x"7d",
          1016 => x"57",
          1017 => x"73",
          1018 => x"ff",
          1019 => x"52",
          1020 => x"fb",
          1021 => x"06",
          1022 => x"2e",
          1023 => x"ff",
          1024 => x"52",
          1025 => x"51",
          1026 => x"74",
          1027 => x"7a",
          1028 => x"f1",
          1029 => x"39",
          1030 => x"98",
          1031 => x"2c",
          1032 => x"b7",
          1033 => x"ab",
          1034 => x"3f",
          1035 => x"52",
          1036 => x"bb",
          1037 => x"39",
          1038 => x"51",
          1039 => x"84",
          1040 => x"83",
          1041 => x"78",
          1042 => x"2b",
          1043 => x"f3",
          1044 => x"07",
          1045 => x"83",
          1046 => x"52",
          1047 => x"99",
          1048 => x"0d",
          1049 => x"08",
          1050 => x"74",
          1051 => x"3f",
          1052 => x"04",
          1053 => x"78",
          1054 => x"84",
          1055 => x"85",
          1056 => x"81",
          1057 => x"70",
          1058 => x"56",
          1059 => x"ff",
          1060 => x"2e",
          1061 => x"80",
          1062 => x"70",
          1063 => x"33",
          1064 => x"2e",
          1065 => x"d4",
          1066 => x"72",
          1067 => x"08",
          1068 => x"84",
          1069 => x"80",
          1070 => x"ff",
          1071 => x"81",
          1072 => x"53",
          1073 => x"88",
          1074 => x"c8",
          1075 => x"39",
          1076 => x"08",
          1077 => x"c8",
          1078 => x"51",
          1079 => x"55",
          1080 => x"b8",
          1081 => x"2e",
          1082 => x"57",
          1083 => x"84",
          1084 => x"88",
          1085 => x"fa",
          1086 => x"7a",
          1087 => x"0b",
          1088 => x"70",
          1089 => x"32",
          1090 => x"51",
          1091 => x"ff",
          1092 => x"2e",
          1093 => x"92",
          1094 => x"81",
          1095 => x"53",
          1096 => x"09",
          1097 => x"38",
          1098 => x"84",
          1099 => x"88",
          1100 => x"73",
          1101 => x"55",
          1102 => x"80",
          1103 => x"74",
          1104 => x"90",
          1105 => x"72",
          1106 => x"e4",
          1107 => x"e3",
          1108 => x"70",
          1109 => x"33",
          1110 => x"e3",
          1111 => x"ff",
          1112 => x"d4",
          1113 => x"73",
          1114 => x"83",
          1115 => x"fa",
          1116 => x"7a",
          1117 => x"70",
          1118 => x"32",
          1119 => x"56",
          1120 => x"56",
          1121 => x"73",
          1122 => x"06",
          1123 => x"2e",
          1124 => x"15",
          1125 => x"88",
          1126 => x"91",
          1127 => x"56",
          1128 => x"74",
          1129 => x"75",
          1130 => x"08",
          1131 => x"8c",
          1132 => x"56",
          1133 => x"e4",
          1134 => x"0d",
          1135 => x"76",
          1136 => x"51",
          1137 => x"54",
          1138 => x"56",
          1139 => x"08",
          1140 => x"15",
          1141 => x"8c",
          1142 => x"56",
          1143 => x"3d",
          1144 => x"11",
          1145 => x"ff",
          1146 => x"32",
          1147 => x"55",
          1148 => x"54",
          1149 => x"72",
          1150 => x"06",
          1151 => x"38",
          1152 => x"81",
          1153 => x"80",
          1154 => x"38",
          1155 => x"33",
          1156 => x"80",
          1157 => x"38",
          1158 => x"0c",
          1159 => x"81",
          1160 => x"0c",
          1161 => x"06",
          1162 => x"b8",
          1163 => x"3d",
          1164 => x"ff",
          1165 => x"72",
          1166 => x"8c",
          1167 => x"05",
          1168 => x"84",
          1169 => x"b8",
          1170 => x"3d",
          1171 => x"51",
          1172 => x"55",
          1173 => x"b8",
          1174 => x"84",
          1175 => x"80",
          1176 => x"38",
          1177 => x"70",
          1178 => x"52",
          1179 => x"08",
          1180 => x"38",
          1181 => x"53",
          1182 => x"34",
          1183 => x"84",
          1184 => x"87",
          1185 => x"74",
          1186 => x"72",
          1187 => x"ff",
          1188 => x"fd",
          1189 => x"77",
          1190 => x"54",
          1191 => x"05",
          1192 => x"70",
          1193 => x"12",
          1194 => x"81",
          1195 => x"51",
          1196 => x"81",
          1197 => x"70",
          1198 => x"84",
          1199 => x"85",
          1200 => x"fc",
          1201 => x"79",
          1202 => x"55",
          1203 => x"80",
          1204 => x"73",
          1205 => x"38",
          1206 => x"93",
          1207 => x"81",
          1208 => x"73",
          1209 => x"55",
          1210 => x"51",
          1211 => x"73",
          1212 => x"0c",
          1213 => x"04",
          1214 => x"73",
          1215 => x"38",
          1216 => x"53",
          1217 => x"ff",
          1218 => x"71",
          1219 => x"ff",
          1220 => x"80",
          1221 => x"ff",
          1222 => x"53",
          1223 => x"73",
          1224 => x"51",
          1225 => x"c7",
          1226 => x"0d",
          1227 => x"53",
          1228 => x"05",
          1229 => x"70",
          1230 => x"12",
          1231 => x"84",
          1232 => x"51",
          1233 => x"04",
          1234 => x"75",
          1235 => x"54",
          1236 => x"81",
          1237 => x"51",
          1238 => x"81",
          1239 => x"70",
          1240 => x"84",
          1241 => x"85",
          1242 => x"fd",
          1243 => x"78",
          1244 => x"55",
          1245 => x"80",
          1246 => x"71",
          1247 => x"53",
          1248 => x"81",
          1249 => x"ff",
          1250 => x"ef",
          1251 => x"b8",
          1252 => x"3d",
          1253 => x"3d",
          1254 => x"7a",
          1255 => x"72",
          1256 => x"38",
          1257 => x"70",
          1258 => x"33",
          1259 => x"71",
          1260 => x"06",
          1261 => x"14",
          1262 => x"2e",
          1263 => x"13",
          1264 => x"38",
          1265 => x"84",
          1266 => x"86",
          1267 => x"72",
          1268 => x"38",
          1269 => x"ff",
          1270 => x"2e",
          1271 => x"15",
          1272 => x"51",
          1273 => x"de",
          1274 => x"31",
          1275 => x"0c",
          1276 => x"04",
          1277 => x"e4",
          1278 => x"0d",
          1279 => x"0d",
          1280 => x"70",
          1281 => x"c1",
          1282 => x"e4",
          1283 => x"e4",
          1284 => x"52",
          1285 => x"d9",
          1286 => x"e4",
          1287 => x"b8",
          1288 => x"2e",
          1289 => x"b8",
          1290 => x"54",
          1291 => x"74",
          1292 => x"84",
          1293 => x"51",
          1294 => x"84",
          1295 => x"54",
          1296 => x"e4",
          1297 => x"0d",
          1298 => x"0d",
          1299 => x"71",
          1300 => x"54",
          1301 => x"9f",
          1302 => x"81",
          1303 => x"51",
          1304 => x"8c",
          1305 => x"52",
          1306 => x"09",
          1307 => x"38",
          1308 => x"75",
          1309 => x"70",
          1310 => x"0c",
          1311 => x"04",
          1312 => x"75",
          1313 => x"55",
          1314 => x"70",
          1315 => x"38",
          1316 => x"81",
          1317 => x"ff",
          1318 => x"f4",
          1319 => x"b8",
          1320 => x"3d",
          1321 => x"3d",
          1322 => x"58",
          1323 => x"76",
          1324 => x"38",
          1325 => x"f5",
          1326 => x"e4",
          1327 => x"12",
          1328 => x"2e",
          1329 => x"51",
          1330 => x"71",
          1331 => x"08",
          1332 => x"52",
          1333 => x"80",
          1334 => x"52",
          1335 => x"80",
          1336 => x"13",
          1337 => x"a0",
          1338 => x"71",
          1339 => x"54",
          1340 => x"74",
          1341 => x"38",
          1342 => x"9f",
          1343 => x"10",
          1344 => x"72",
          1345 => x"9f",
          1346 => x"06",
          1347 => x"75",
          1348 => x"1c",
          1349 => x"52",
          1350 => x"53",
          1351 => x"73",
          1352 => x"52",
          1353 => x"e4",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"80",
          1357 => x"30",
          1358 => x"80",
          1359 => x"2b",
          1360 => x"75",
          1361 => x"83",
          1362 => x"70",
          1363 => x"25",
          1364 => x"71",
          1365 => x"2a",
          1366 => x"06",
          1367 => x"80",
          1368 => x"84",
          1369 => x"71",
          1370 => x"75",
          1371 => x"8c",
          1372 => x"70",
          1373 => x"82",
          1374 => x"71",
          1375 => x"2a",
          1376 => x"81",
          1377 => x"82",
          1378 => x"75",
          1379 => x"b8",
          1380 => x"52",
          1381 => x"54",
          1382 => x"55",
          1383 => x"56",
          1384 => x"51",
          1385 => x"52",
          1386 => x"04",
          1387 => x"75",
          1388 => x"71",
          1389 => x"81",
          1390 => x"b8",
          1391 => x"29",
          1392 => x"84",
          1393 => x"53",
          1394 => x"04",
          1395 => x"78",
          1396 => x"a0",
          1397 => x"2e",
          1398 => x"51",
          1399 => x"84",
          1400 => x"53",
          1401 => x"73",
          1402 => x"38",
          1403 => x"bd",
          1404 => x"b8",
          1405 => x"52",
          1406 => x"9f",
          1407 => x"38",
          1408 => x"9f",
          1409 => x"81",
          1410 => x"2a",
          1411 => x"76",
          1412 => x"54",
          1413 => x"56",
          1414 => x"a8",
          1415 => x"74",
          1416 => x"74",
          1417 => x"78",
          1418 => x"11",
          1419 => x"81",
          1420 => x"06",
          1421 => x"ff",
          1422 => x"52",
          1423 => x"55",
          1424 => x"38",
          1425 => x"e4",
          1426 => x"0d",
          1427 => x"0d",
          1428 => x"7a",
          1429 => x"9f",
          1430 => x"7c",
          1431 => x"32",
          1432 => x"71",
          1433 => x"72",
          1434 => x"59",
          1435 => x"56",
          1436 => x"84",
          1437 => x"75",
          1438 => x"84",
          1439 => x"88",
          1440 => x"f7",
          1441 => x"7d",
          1442 => x"70",
          1443 => x"08",
          1444 => x"56",
          1445 => x"2e",
          1446 => x"8f",
          1447 => x"70",
          1448 => x"33",
          1449 => x"a0",
          1450 => x"73",
          1451 => x"f5",
          1452 => x"2e",
          1453 => x"d0",
          1454 => x"56",
          1455 => x"80",
          1456 => x"58",
          1457 => x"74",
          1458 => x"38",
          1459 => x"27",
          1460 => x"14",
          1461 => x"06",
          1462 => x"14",
          1463 => x"06",
          1464 => x"73",
          1465 => x"f9",
          1466 => x"ff",
          1467 => x"89",
          1468 => x"89",
          1469 => x"27",
          1470 => x"77",
          1471 => x"81",
          1472 => x"0c",
          1473 => x"56",
          1474 => x"26",
          1475 => x"78",
          1476 => x"38",
          1477 => x"75",
          1478 => x"56",
          1479 => x"e4",
          1480 => x"0d",
          1481 => x"16",
          1482 => x"70",
          1483 => x"59",
          1484 => x"09",
          1485 => x"ff",
          1486 => x"70",
          1487 => x"33",
          1488 => x"80",
          1489 => x"38",
          1490 => x"80",
          1491 => x"38",
          1492 => x"74",
          1493 => x"d0",
          1494 => x"56",
          1495 => x"73",
          1496 => x"38",
          1497 => x"e4",
          1498 => x"0d",
          1499 => x"81",
          1500 => x"0c",
          1501 => x"55",
          1502 => x"ca",
          1503 => x"84",
          1504 => x"8b",
          1505 => x"f7",
          1506 => x"7d",
          1507 => x"70",
          1508 => x"08",
          1509 => x"56",
          1510 => x"2e",
          1511 => x"8f",
          1512 => x"70",
          1513 => x"33",
          1514 => x"a0",
          1515 => x"73",
          1516 => x"f5",
          1517 => x"2e",
          1518 => x"d0",
          1519 => x"56",
          1520 => x"80",
          1521 => x"58",
          1522 => x"74",
          1523 => x"38",
          1524 => x"27",
          1525 => x"14",
          1526 => x"06",
          1527 => x"14",
          1528 => x"06",
          1529 => x"73",
          1530 => x"f9",
          1531 => x"ff",
          1532 => x"89",
          1533 => x"89",
          1534 => x"27",
          1535 => x"77",
          1536 => x"81",
          1537 => x"0c",
          1538 => x"56",
          1539 => x"26",
          1540 => x"78",
          1541 => x"38",
          1542 => x"75",
          1543 => x"56",
          1544 => x"e4",
          1545 => x"0d",
          1546 => x"16",
          1547 => x"70",
          1548 => x"59",
          1549 => x"09",
          1550 => x"ff",
          1551 => x"70",
          1552 => x"33",
          1553 => x"80",
          1554 => x"38",
          1555 => x"80",
          1556 => x"38",
          1557 => x"74",
          1558 => x"d0",
          1559 => x"56",
          1560 => x"73",
          1561 => x"38",
          1562 => x"e4",
          1563 => x"0d",
          1564 => x"81",
          1565 => x"0c",
          1566 => x"55",
          1567 => x"ca",
          1568 => x"84",
          1569 => x"8b",
          1570 => x"80",
          1571 => x"84",
          1572 => x"81",
          1573 => x"b8",
          1574 => x"ff",
          1575 => x"52",
          1576 => x"8c",
          1577 => x"10",
          1578 => x"05",
          1579 => x"04",
          1580 => x"51",
          1581 => x"83",
          1582 => x"83",
          1583 => x"ef",
          1584 => x"3d",
          1585 => x"ce",
          1586 => x"a8",
          1587 => x"0d",
          1588 => x"cc",
          1589 => x"3f",
          1590 => x"04",
          1591 => x"51",
          1592 => x"83",
          1593 => x"83",
          1594 => x"ef",
          1595 => x"3d",
          1596 => x"cf",
          1597 => x"fc",
          1598 => x"0d",
          1599 => x"a4",
          1600 => x"3f",
          1601 => x"04",
          1602 => x"51",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ee",
          1606 => x"3d",
          1607 => x"cf",
          1608 => x"d0",
          1609 => x"0d",
          1610 => x"94",
          1611 => x"3f",
          1612 => x"04",
          1613 => x"51",
          1614 => x"83",
          1615 => x"83",
          1616 => x"ee",
          1617 => x"3d",
          1618 => x"d0",
          1619 => x"a4",
          1620 => x"0d",
          1621 => x"e8",
          1622 => x"3f",
          1623 => x"04",
          1624 => x"51",
          1625 => x"83",
          1626 => x"83",
          1627 => x"ee",
          1628 => x"3d",
          1629 => x"d1",
          1630 => x"f8",
          1631 => x"0d",
          1632 => x"a8",
          1633 => x"3f",
          1634 => x"04",
          1635 => x"51",
          1636 => x"83",
          1637 => x"ec",
          1638 => x"02",
          1639 => x"e3",
          1640 => x"58",
          1641 => x"30",
          1642 => x"73",
          1643 => x"57",
          1644 => x"75",
          1645 => x"83",
          1646 => x"74",
          1647 => x"81",
          1648 => x"55",
          1649 => x"80",
          1650 => x"53",
          1651 => x"3d",
          1652 => x"82",
          1653 => x"84",
          1654 => x"57",
          1655 => x"08",
          1656 => x"d0",
          1657 => x"82",
          1658 => x"76",
          1659 => x"07",
          1660 => x"30",
          1661 => x"72",
          1662 => x"57",
          1663 => x"2e",
          1664 => x"c0",
          1665 => x"55",
          1666 => x"26",
          1667 => x"74",
          1668 => x"e8",
          1669 => x"8e",
          1670 => x"e4",
          1671 => x"d1",
          1672 => x"52",
          1673 => x"51",
          1674 => x"76",
          1675 => x"0c",
          1676 => x"04",
          1677 => x"08",
          1678 => x"88",
          1679 => x"e4",
          1680 => x"3d",
          1681 => x"84",
          1682 => x"52",
          1683 => x"9d",
          1684 => x"b8",
          1685 => x"84",
          1686 => x"ff",
          1687 => x"55",
          1688 => x"ff",
          1689 => x"19",
          1690 => x"59",
          1691 => x"e8",
          1692 => x"f4",
          1693 => x"b8",
          1694 => x"78",
          1695 => x"3f",
          1696 => x"08",
          1697 => x"e4",
          1698 => x"83",
          1699 => x"de",
          1700 => x"97",
          1701 => x"0d",
          1702 => x"05",
          1703 => x"58",
          1704 => x"80",
          1705 => x"7a",
          1706 => x"3f",
          1707 => x"08",
          1708 => x"80",
          1709 => x"76",
          1710 => x"38",
          1711 => x"e4",
          1712 => x"0d",
          1713 => x"84",
          1714 => x"61",
          1715 => x"84",
          1716 => x"7f",
          1717 => x"78",
          1718 => x"e4",
          1719 => x"e4",
          1720 => x"0d",
          1721 => x"0d",
          1722 => x"02",
          1723 => x"cf",
          1724 => x"73",
          1725 => x"5f",
          1726 => x"5d",
          1727 => x"2e",
          1728 => x"7a",
          1729 => x"ec",
          1730 => x"3f",
          1731 => x"51",
          1732 => x"80",
          1733 => x"27",
          1734 => x"90",
          1735 => x"38",
          1736 => x"82",
          1737 => x"18",
          1738 => x"27",
          1739 => x"72",
          1740 => x"d1",
          1741 => x"d1",
          1742 => x"84",
          1743 => x"53",
          1744 => x"ec",
          1745 => x"74",
          1746 => x"83",
          1747 => x"dd",
          1748 => x"56",
          1749 => x"80",
          1750 => x"18",
          1751 => x"53",
          1752 => x"7a",
          1753 => x"81",
          1754 => x"9f",
          1755 => x"38",
          1756 => x"73",
          1757 => x"ff",
          1758 => x"74",
          1759 => x"38",
          1760 => x"27",
          1761 => x"84",
          1762 => x"52",
          1763 => x"df",
          1764 => x"56",
          1765 => x"c2",
          1766 => x"84",
          1767 => x"3f",
          1768 => x"1c",
          1769 => x"51",
          1770 => x"84",
          1771 => x"98",
          1772 => x"2c",
          1773 => x"a0",
          1774 => x"38",
          1775 => x"82",
          1776 => x"1e",
          1777 => x"26",
          1778 => x"ff",
          1779 => x"e4",
          1780 => x"0d",
          1781 => x"88",
          1782 => x"3f",
          1783 => x"d4",
          1784 => x"54",
          1785 => x"87",
          1786 => x"26",
          1787 => x"fe",
          1788 => x"d2",
          1789 => x"91",
          1790 => x"84",
          1791 => x"53",
          1792 => x"ea",
          1793 => x"79",
          1794 => x"38",
          1795 => x"72",
          1796 => x"38",
          1797 => x"83",
          1798 => x"db",
          1799 => x"14",
          1800 => x"08",
          1801 => x"51",
          1802 => x"78",
          1803 => x"38",
          1804 => x"83",
          1805 => x"db",
          1806 => x"14",
          1807 => x"08",
          1808 => x"51",
          1809 => x"73",
          1810 => x"ff",
          1811 => x"53",
          1812 => x"df",
          1813 => x"52",
          1814 => x"51",
          1815 => x"84",
          1816 => x"c8",
          1817 => x"a0",
          1818 => x"3f",
          1819 => x"dd",
          1820 => x"39",
          1821 => x"08",
          1822 => x"e9",
          1823 => x"16",
          1824 => x"39",
          1825 => x"3f",
          1826 => x"08",
          1827 => x"53",
          1828 => x"a8",
          1829 => x"38",
          1830 => x"80",
          1831 => x"81",
          1832 => x"38",
          1833 => x"db",
          1834 => x"9b",
          1835 => x"b8",
          1836 => x"2b",
          1837 => x"70",
          1838 => x"30",
          1839 => x"70",
          1840 => x"07",
          1841 => x"06",
          1842 => x"59",
          1843 => x"72",
          1844 => x"e8",
          1845 => x"9a",
          1846 => x"b8",
          1847 => x"2b",
          1848 => x"70",
          1849 => x"30",
          1850 => x"70",
          1851 => x"07",
          1852 => x"06",
          1853 => x"59",
          1854 => x"80",
          1855 => x"a9",
          1856 => x"39",
          1857 => x"b8",
          1858 => x"3d",
          1859 => x"3d",
          1860 => x"96",
          1861 => x"aa",
          1862 => x"51",
          1863 => x"83",
          1864 => x"9c",
          1865 => x"51",
          1866 => x"72",
          1867 => x"81",
          1868 => x"71",
          1869 => x"72",
          1870 => x"81",
          1871 => x"71",
          1872 => x"72",
          1873 => x"81",
          1874 => x"71",
          1875 => x"72",
          1876 => x"81",
          1877 => x"71",
          1878 => x"72",
          1879 => x"81",
          1880 => x"71",
          1881 => x"72",
          1882 => x"81",
          1883 => x"71",
          1884 => x"72",
          1885 => x"81",
          1886 => x"71",
          1887 => x"88",
          1888 => x"53",
          1889 => x"a9",
          1890 => x"3d",
          1891 => x"51",
          1892 => x"83",
          1893 => x"9c",
          1894 => x"51",
          1895 => x"a9",
          1896 => x"3d",
          1897 => x"51",
          1898 => x"83",
          1899 => x"9b",
          1900 => x"51",
          1901 => x"72",
          1902 => x"06",
          1903 => x"2e",
          1904 => x"39",
          1905 => x"c3",
          1906 => x"9c",
          1907 => x"3f",
          1908 => x"b7",
          1909 => x"2a",
          1910 => x"51",
          1911 => x"2e",
          1912 => x"c2",
          1913 => x"9b",
          1914 => x"d3",
          1915 => x"b3",
          1916 => x"9b",
          1917 => x"86",
          1918 => x"06",
          1919 => x"80",
          1920 => x"38",
          1921 => x"81",
          1922 => x"3f",
          1923 => x"51",
          1924 => x"80",
          1925 => x"3f",
          1926 => x"70",
          1927 => x"52",
          1928 => x"fe",
          1929 => x"bd",
          1930 => x"9a",
          1931 => x"d3",
          1932 => x"ef",
          1933 => x"9a",
          1934 => x"84",
          1935 => x"06",
          1936 => x"80",
          1937 => x"38",
          1938 => x"81",
          1939 => x"3f",
          1940 => x"51",
          1941 => x"80",
          1942 => x"3f",
          1943 => x"70",
          1944 => x"52",
          1945 => x"fd",
          1946 => x"bd",
          1947 => x"9a",
          1948 => x"d3",
          1949 => x"ab",
          1950 => x"9a",
          1951 => x"82",
          1952 => x"06",
          1953 => x"80",
          1954 => x"38",
          1955 => x"ca",
          1956 => x"70",
          1957 => x"61",
          1958 => x"0c",
          1959 => x"60",
          1960 => x"fb",
          1961 => x"e4",
          1962 => x"06",
          1963 => x"59",
          1964 => x"84",
          1965 => x"d4",
          1966 => x"b8",
          1967 => x"43",
          1968 => x"51",
          1969 => x"7e",
          1970 => x"53",
          1971 => x"51",
          1972 => x"0b",
          1973 => x"d8",
          1974 => x"ff",
          1975 => x"79",
          1976 => x"f1",
          1977 => x"2e",
          1978 => x"78",
          1979 => x"5e",
          1980 => x"83",
          1981 => x"70",
          1982 => x"80",
          1983 => x"38",
          1984 => x"7b",
          1985 => x"81",
          1986 => x"81",
          1987 => x"5d",
          1988 => x"2e",
          1989 => x"5c",
          1990 => x"be",
          1991 => x"29",
          1992 => x"05",
          1993 => x"5b",
          1994 => x"84",
          1995 => x"84",
          1996 => x"54",
          1997 => x"08",
          1998 => x"da",
          1999 => x"e4",
          2000 => x"84",
          2001 => x"7d",
          2002 => x"80",
          2003 => x"70",
          2004 => x"5d",
          2005 => x"27",
          2006 => x"3d",
          2007 => x"80",
          2008 => x"38",
          2009 => x"7e",
          2010 => x"3f",
          2011 => x"08",
          2012 => x"e4",
          2013 => x"8d",
          2014 => x"b8",
          2015 => x"b8",
          2016 => x"05",
          2017 => x"3f",
          2018 => x"08",
          2019 => x"5c",
          2020 => x"2e",
          2021 => x"84",
          2022 => x"51",
          2023 => x"84",
          2024 => x"8f",
          2025 => x"38",
          2026 => x"3d",
          2027 => x"82",
          2028 => x"38",
          2029 => x"8c",
          2030 => x"81",
          2031 => x"38",
          2032 => x"53",
          2033 => x"52",
          2034 => x"dd",
          2035 => x"a0",
          2036 => x"94",
          2037 => x"67",
          2038 => x"90",
          2039 => x"90",
          2040 => x"7c",
          2041 => x"3f",
          2042 => x"08",
          2043 => x"08",
          2044 => x"70",
          2045 => x"25",
          2046 => x"42",
          2047 => x"83",
          2048 => x"81",
          2049 => x"06",
          2050 => x"2e",
          2051 => x"1b",
          2052 => x"06",
          2053 => x"ff",
          2054 => x"81",
          2055 => x"32",
          2056 => x"81",
          2057 => x"ff",
          2058 => x"38",
          2059 => x"94",
          2060 => x"d5",
          2061 => x"d1",
          2062 => x"80",
          2063 => x"52",
          2064 => x"bc",
          2065 => x"83",
          2066 => x"70",
          2067 => x"5b",
          2068 => x"91",
          2069 => x"83",
          2070 => x"84",
          2071 => x"82",
          2072 => x"84",
          2073 => x"80",
          2074 => x"0b",
          2075 => x"ed",
          2076 => x"cf",
          2077 => x"f8",
          2078 => x"82",
          2079 => x"84",
          2080 => x"80",
          2081 => x"84",
          2082 => x"51",
          2083 => x"0b",
          2084 => x"d8",
          2085 => x"ff",
          2086 => x"7d",
          2087 => x"81",
          2088 => x"38",
          2089 => x"cf",
          2090 => x"a1",
          2091 => x"0b",
          2092 => x"ed",
          2093 => x"d4",
          2094 => x"f8",
          2095 => x"a7",
          2096 => x"70",
          2097 => x"fc",
          2098 => x"39",
          2099 => x"0c",
          2100 => x"59",
          2101 => x"26",
          2102 => x"78",
          2103 => x"be",
          2104 => x"79",
          2105 => x"53",
          2106 => x"52",
          2107 => x"fb",
          2108 => x"7e",
          2109 => x"90",
          2110 => x"f3",
          2111 => x"e4",
          2112 => x"09",
          2113 => x"ae",
          2114 => x"9a",
          2115 => x"41",
          2116 => x"83",
          2117 => x"de",
          2118 => x"51",
          2119 => x"3f",
          2120 => x"83",
          2121 => x"7b",
          2122 => x"ac",
          2123 => x"83",
          2124 => x"7c",
          2125 => x"3f",
          2126 => x"81",
          2127 => x"fa",
          2128 => x"dd",
          2129 => x"39",
          2130 => x"51",
          2131 => x"fa",
          2132 => x"8d",
          2133 => x"e8",
          2134 => x"c0",
          2135 => x"3f",
          2136 => x"04",
          2137 => x"51",
          2138 => x"d0",
          2139 => x"d0",
          2140 => x"ff",
          2141 => x"ff",
          2142 => x"ec",
          2143 => x"b8",
          2144 => x"2e",
          2145 => x"68",
          2146 => x"f0",
          2147 => x"3f",
          2148 => x"2d",
          2149 => x"08",
          2150 => x"a4",
          2151 => x"e4",
          2152 => x"d6",
          2153 => x"e1",
          2154 => x"39",
          2155 => x"84",
          2156 => x"80",
          2157 => x"cf",
          2158 => x"e4",
          2159 => x"f9",
          2160 => x"52",
          2161 => x"51",
          2162 => x"68",
          2163 => x"b8",
          2164 => x"11",
          2165 => x"05",
          2166 => x"3f",
          2167 => x"08",
          2168 => x"dc",
          2169 => x"fe",
          2170 => x"ff",
          2171 => x"e9",
          2172 => x"b8",
          2173 => x"d0",
          2174 => x"78",
          2175 => x"52",
          2176 => x"51",
          2177 => x"84",
          2178 => x"53",
          2179 => x"7e",
          2180 => x"3f",
          2181 => x"33",
          2182 => x"2e",
          2183 => x"78",
          2184 => x"d3",
          2185 => x"05",
          2186 => x"cf",
          2187 => x"fe",
          2188 => x"ff",
          2189 => x"e8",
          2190 => x"b8",
          2191 => x"2e",
          2192 => x"b8",
          2193 => x"11",
          2194 => x"05",
          2195 => x"3f",
          2196 => x"08",
          2197 => x"64",
          2198 => x"53",
          2199 => x"d6",
          2200 => x"a5",
          2201 => x"c4",
          2202 => x"f8",
          2203 => x"cf",
          2204 => x"48",
          2205 => x"78",
          2206 => x"c4",
          2207 => x"26",
          2208 => x"64",
          2209 => x"46",
          2210 => x"b8",
          2211 => x"11",
          2212 => x"05",
          2213 => x"3f",
          2214 => x"08",
          2215 => x"a0",
          2216 => x"fe",
          2217 => x"ff",
          2218 => x"e9",
          2219 => x"b8",
          2220 => x"2e",
          2221 => x"b8",
          2222 => x"11",
          2223 => x"05",
          2224 => x"3f",
          2225 => x"08",
          2226 => x"f4",
          2227 => x"e0",
          2228 => x"3f",
          2229 => x"59",
          2230 => x"83",
          2231 => x"70",
          2232 => x"5f",
          2233 => x"7d",
          2234 => x"7a",
          2235 => x"78",
          2236 => x"52",
          2237 => x"51",
          2238 => x"66",
          2239 => x"81",
          2240 => x"47",
          2241 => x"b8",
          2242 => x"11",
          2243 => x"05",
          2244 => x"3f",
          2245 => x"08",
          2246 => x"a4",
          2247 => x"fe",
          2248 => x"ff",
          2249 => x"e8",
          2250 => x"b8",
          2251 => x"2e",
          2252 => x"b8",
          2253 => x"11",
          2254 => x"05",
          2255 => x"3f",
          2256 => x"08",
          2257 => x"f8",
          2258 => x"8c",
          2259 => x"3f",
          2260 => x"67",
          2261 => x"38",
          2262 => x"70",
          2263 => x"33",
          2264 => x"81",
          2265 => x"39",
          2266 => x"84",
          2267 => x"80",
          2268 => x"93",
          2269 => x"e4",
          2270 => x"f6",
          2271 => x"3d",
          2272 => x"53",
          2273 => x"51",
          2274 => x"84",
          2275 => x"b1",
          2276 => x"33",
          2277 => x"d7",
          2278 => x"ed",
          2279 => x"c4",
          2280 => x"f8",
          2281 => x"cc",
          2282 => x"48",
          2283 => x"78",
          2284 => x"8c",
          2285 => x"26",
          2286 => x"68",
          2287 => x"d1",
          2288 => x"02",
          2289 => x"33",
          2290 => x"81",
          2291 => x"3d",
          2292 => x"53",
          2293 => x"51",
          2294 => x"84",
          2295 => x"80",
          2296 => x"38",
          2297 => x"80",
          2298 => x"79",
          2299 => x"05",
          2300 => x"fe",
          2301 => x"ff",
          2302 => x"e7",
          2303 => x"b8",
          2304 => x"bd",
          2305 => x"39",
          2306 => x"84",
          2307 => x"80",
          2308 => x"f3",
          2309 => x"e4",
          2310 => x"f5",
          2311 => x"3d",
          2312 => x"53",
          2313 => x"51",
          2314 => x"84",
          2315 => x"80",
          2316 => x"38",
          2317 => x"f8",
          2318 => x"80",
          2319 => x"c7",
          2320 => x"e4",
          2321 => x"84",
          2322 => x"46",
          2323 => x"51",
          2324 => x"68",
          2325 => x"78",
          2326 => x"38",
          2327 => x"79",
          2328 => x"5b",
          2329 => x"26",
          2330 => x"51",
          2331 => x"f4",
          2332 => x"3d",
          2333 => x"51",
          2334 => x"84",
          2335 => x"b9",
          2336 => x"05",
          2337 => x"d8",
          2338 => x"84",
          2339 => x"52",
          2340 => x"83",
          2341 => x"e4",
          2342 => x"f4",
          2343 => x"b8",
          2344 => x"e7",
          2345 => x"98",
          2346 => x"ff",
          2347 => x"ff",
          2348 => x"e5",
          2349 => x"b8",
          2350 => x"38",
          2351 => x"33",
          2352 => x"2e",
          2353 => x"83",
          2354 => x"49",
          2355 => x"fc",
          2356 => x"80",
          2357 => x"af",
          2358 => x"e4",
          2359 => x"83",
          2360 => x"5a",
          2361 => x"83",
          2362 => x"f1",
          2363 => x"b8",
          2364 => x"11",
          2365 => x"05",
          2366 => x"3f",
          2367 => x"08",
          2368 => x"38",
          2369 => x"5c",
          2370 => x"83",
          2371 => x"7a",
          2372 => x"30",
          2373 => x"9f",
          2374 => x"5c",
          2375 => x"80",
          2376 => x"7a",
          2377 => x"38",
          2378 => x"d7",
          2379 => x"c4",
          2380 => x"68",
          2381 => x"66",
          2382 => x"eb",
          2383 => x"d7",
          2384 => x"b0",
          2385 => x"39",
          2386 => x"0c",
          2387 => x"05",
          2388 => x"fe",
          2389 => x"ff",
          2390 => x"e2",
          2391 => x"b8",
          2392 => x"2e",
          2393 => x"64",
          2394 => x"59",
          2395 => x"45",
          2396 => x"f0",
          2397 => x"80",
          2398 => x"87",
          2399 => x"e4",
          2400 => x"f2",
          2401 => x"5e",
          2402 => x"05",
          2403 => x"82",
          2404 => x"7d",
          2405 => x"fe",
          2406 => x"ff",
          2407 => x"e1",
          2408 => x"b8",
          2409 => x"2e",
          2410 => x"64",
          2411 => x"ce",
          2412 => x"70",
          2413 => x"23",
          2414 => x"3d",
          2415 => x"53",
          2416 => x"51",
          2417 => x"84",
          2418 => x"ff",
          2419 => x"f0",
          2420 => x"fe",
          2421 => x"ff",
          2422 => x"e3",
          2423 => x"b8",
          2424 => x"2e",
          2425 => x"68",
          2426 => x"db",
          2427 => x"34",
          2428 => x"49",
          2429 => x"b8",
          2430 => x"11",
          2431 => x"05",
          2432 => x"3f",
          2433 => x"08",
          2434 => x"98",
          2435 => x"71",
          2436 => x"84",
          2437 => x"59",
          2438 => x"7a",
          2439 => x"81",
          2440 => x"38",
          2441 => x"d5",
          2442 => x"53",
          2443 => x"52",
          2444 => x"f5",
          2445 => x"39",
          2446 => x"51",
          2447 => x"f3",
          2448 => x"d7",
          2449 => x"ac",
          2450 => x"39",
          2451 => x"f0",
          2452 => x"80",
          2453 => x"ab",
          2454 => x"e4",
          2455 => x"b8",
          2456 => x"02",
          2457 => x"22",
          2458 => x"05",
          2459 => x"45",
          2460 => x"83",
          2461 => x"5c",
          2462 => x"80",
          2463 => x"f1",
          2464 => x"fc",
          2465 => x"f1",
          2466 => x"7b",
          2467 => x"38",
          2468 => x"08",
          2469 => x"39",
          2470 => x"51",
          2471 => x"64",
          2472 => x"39",
          2473 => x"51",
          2474 => x"64",
          2475 => x"39",
          2476 => x"33",
          2477 => x"2e",
          2478 => x"f1",
          2479 => x"fc",
          2480 => x"d8",
          2481 => x"ac",
          2482 => x"39",
          2483 => x"33",
          2484 => x"2e",
          2485 => x"f1",
          2486 => x"fc",
          2487 => x"f1",
          2488 => x"7d",
          2489 => x"38",
          2490 => x"08",
          2491 => x"39",
          2492 => x"33",
          2493 => x"2e",
          2494 => x"f1",
          2495 => x"fb",
          2496 => x"f1",
          2497 => x"7c",
          2498 => x"38",
          2499 => x"08",
          2500 => x"39",
          2501 => x"33",
          2502 => x"2e",
          2503 => x"f1",
          2504 => x"fb",
          2505 => x"f1",
          2506 => x"80",
          2507 => x"9c",
          2508 => x"d0",
          2509 => x"47",
          2510 => x"f3",
          2511 => x"0b",
          2512 => x"34",
          2513 => x"8c",
          2514 => x"57",
          2515 => x"52",
          2516 => x"d2",
          2517 => x"e4",
          2518 => x"77",
          2519 => x"87",
          2520 => x"75",
          2521 => x"3f",
          2522 => x"e4",
          2523 => x"0c",
          2524 => x"9c",
          2525 => x"57",
          2526 => x"52",
          2527 => x"a6",
          2528 => x"e4",
          2529 => x"77",
          2530 => x"87",
          2531 => x"75",
          2532 => x"3f",
          2533 => x"e4",
          2534 => x"0c",
          2535 => x"0b",
          2536 => x"84",
          2537 => x"83",
          2538 => x"94",
          2539 => x"bc",
          2540 => x"c7",
          2541 => x"02",
          2542 => x"05",
          2543 => x"84",
          2544 => x"89",
          2545 => x"13",
          2546 => x"0c",
          2547 => x"0c",
          2548 => x"3f",
          2549 => x"95",
          2550 => x"8d",
          2551 => x"3f",
          2552 => x"52",
          2553 => x"51",
          2554 => x"83",
          2555 => x"22",
          2556 => x"87",
          2557 => x"ac",
          2558 => x"b8",
          2559 => x"33",
          2560 => x"c0",
          2561 => x"3f",
          2562 => x"ed",
          2563 => x"04",
          2564 => x"77",
          2565 => x"56",
          2566 => x"53",
          2567 => x"81",
          2568 => x"33",
          2569 => x"06",
          2570 => x"a0",
          2571 => x"06",
          2572 => x"15",
          2573 => x"81",
          2574 => x"53",
          2575 => x"2e",
          2576 => x"81",
          2577 => x"73",
          2578 => x"82",
          2579 => x"72",
          2580 => x"e7",
          2581 => x"33",
          2582 => x"06",
          2583 => x"70",
          2584 => x"38",
          2585 => x"80",
          2586 => x"73",
          2587 => x"38",
          2588 => x"e1",
          2589 => x"81",
          2590 => x"54",
          2591 => x"09",
          2592 => x"38",
          2593 => x"a2",
          2594 => x"70",
          2595 => x"07",
          2596 => x"72",
          2597 => x"38",
          2598 => x"81",
          2599 => x"71",
          2600 => x"51",
          2601 => x"e4",
          2602 => x"0d",
          2603 => x"2e",
          2604 => x"80",
          2605 => x"38",
          2606 => x"80",
          2607 => x"81",
          2608 => x"54",
          2609 => x"2e",
          2610 => x"54",
          2611 => x"15",
          2612 => x"53",
          2613 => x"2e",
          2614 => x"fe",
          2615 => x"39",
          2616 => x"76",
          2617 => x"8b",
          2618 => x"84",
          2619 => x"86",
          2620 => x"86",
          2621 => x"52",
          2622 => x"87",
          2623 => x"e4",
          2624 => x"e5",
          2625 => x"b8",
          2626 => x"3d",
          2627 => x"3d",
          2628 => x"11",
          2629 => x"52",
          2630 => x"70",
          2631 => x"98",
          2632 => x"33",
          2633 => x"82",
          2634 => x"26",
          2635 => x"84",
          2636 => x"83",
          2637 => x"26",
          2638 => x"85",
          2639 => x"84",
          2640 => x"26",
          2641 => x"86",
          2642 => x"85",
          2643 => x"26",
          2644 => x"88",
          2645 => x"86",
          2646 => x"e7",
          2647 => x"38",
          2648 => x"54",
          2649 => x"87",
          2650 => x"cc",
          2651 => x"87",
          2652 => x"0c",
          2653 => x"c0",
          2654 => x"82",
          2655 => x"c0",
          2656 => x"83",
          2657 => x"c0",
          2658 => x"84",
          2659 => x"c0",
          2660 => x"85",
          2661 => x"c0",
          2662 => x"86",
          2663 => x"c0",
          2664 => x"74",
          2665 => x"a4",
          2666 => x"c0",
          2667 => x"80",
          2668 => x"98",
          2669 => x"52",
          2670 => x"e4",
          2671 => x"0d",
          2672 => x"0d",
          2673 => x"c0",
          2674 => x"81",
          2675 => x"c0",
          2676 => x"5e",
          2677 => x"87",
          2678 => x"08",
          2679 => x"1c",
          2680 => x"98",
          2681 => x"79",
          2682 => x"87",
          2683 => x"08",
          2684 => x"1c",
          2685 => x"98",
          2686 => x"79",
          2687 => x"87",
          2688 => x"08",
          2689 => x"1c",
          2690 => x"98",
          2691 => x"7b",
          2692 => x"87",
          2693 => x"08",
          2694 => x"1c",
          2695 => x"0c",
          2696 => x"ff",
          2697 => x"83",
          2698 => x"58",
          2699 => x"57",
          2700 => x"56",
          2701 => x"55",
          2702 => x"54",
          2703 => x"53",
          2704 => x"ff",
          2705 => x"d8",
          2706 => x"bf",
          2707 => x"3d",
          2708 => x"3d",
          2709 => x"05",
          2710 => x"81",
          2711 => x"72",
          2712 => x"b0",
          2713 => x"e4",
          2714 => x"70",
          2715 => x"52",
          2716 => x"09",
          2717 => x"38",
          2718 => x"e3",
          2719 => x"b8",
          2720 => x"3d",
          2721 => x"51",
          2722 => x"3f",
          2723 => x"08",
          2724 => x"98",
          2725 => x"71",
          2726 => x"81",
          2727 => x"72",
          2728 => x"f0",
          2729 => x"e4",
          2730 => x"70",
          2731 => x"52",
          2732 => x"d2",
          2733 => x"fd",
          2734 => x"70",
          2735 => x"88",
          2736 => x"51",
          2737 => x"3f",
          2738 => x"08",
          2739 => x"98",
          2740 => x"71",
          2741 => x"38",
          2742 => x"81",
          2743 => x"83",
          2744 => x"38",
          2745 => x"e4",
          2746 => x"0d",
          2747 => x"0d",
          2748 => x"33",
          2749 => x"33",
          2750 => x"06",
          2751 => x"70",
          2752 => x"f4",
          2753 => x"94",
          2754 => x"96",
          2755 => x"06",
          2756 => x"70",
          2757 => x"38",
          2758 => x"70",
          2759 => x"51",
          2760 => x"72",
          2761 => x"06",
          2762 => x"2e",
          2763 => x"93",
          2764 => x"52",
          2765 => x"73",
          2766 => x"51",
          2767 => x"80",
          2768 => x"2e",
          2769 => x"c0",
          2770 => x"74",
          2771 => x"84",
          2772 => x"86",
          2773 => x"71",
          2774 => x"81",
          2775 => x"70",
          2776 => x"81",
          2777 => x"53",
          2778 => x"cb",
          2779 => x"2a",
          2780 => x"71",
          2781 => x"38",
          2782 => x"84",
          2783 => x"2a",
          2784 => x"53",
          2785 => x"cf",
          2786 => x"ff",
          2787 => x"8f",
          2788 => x"30",
          2789 => x"51",
          2790 => x"83",
          2791 => x"83",
          2792 => x"fa",
          2793 => x"55",
          2794 => x"70",
          2795 => x"70",
          2796 => x"e7",
          2797 => x"83",
          2798 => x"70",
          2799 => x"54",
          2800 => x"80",
          2801 => x"38",
          2802 => x"94",
          2803 => x"2a",
          2804 => x"53",
          2805 => x"80",
          2806 => x"71",
          2807 => x"81",
          2808 => x"70",
          2809 => x"81",
          2810 => x"53",
          2811 => x"8a",
          2812 => x"2a",
          2813 => x"71",
          2814 => x"81",
          2815 => x"87",
          2816 => x"52",
          2817 => x"86",
          2818 => x"94",
          2819 => x"72",
          2820 => x"75",
          2821 => x"73",
          2822 => x"76",
          2823 => x"0c",
          2824 => x"04",
          2825 => x"70",
          2826 => x"51",
          2827 => x"72",
          2828 => x"06",
          2829 => x"2e",
          2830 => x"93",
          2831 => x"52",
          2832 => x"ff",
          2833 => x"c0",
          2834 => x"70",
          2835 => x"81",
          2836 => x"52",
          2837 => x"d7",
          2838 => x"0d",
          2839 => x"80",
          2840 => x"2a",
          2841 => x"52",
          2842 => x"84",
          2843 => x"c0",
          2844 => x"83",
          2845 => x"87",
          2846 => x"08",
          2847 => x"0c",
          2848 => x"94",
          2849 => x"a8",
          2850 => x"9e",
          2851 => x"f1",
          2852 => x"c0",
          2853 => x"83",
          2854 => x"87",
          2855 => x"08",
          2856 => x"0c",
          2857 => x"ac",
          2858 => x"b8",
          2859 => x"9e",
          2860 => x"f1",
          2861 => x"c0",
          2862 => x"83",
          2863 => x"87",
          2864 => x"08",
          2865 => x"0c",
          2866 => x"bc",
          2867 => x"c8",
          2868 => x"9e",
          2869 => x"f1",
          2870 => x"c0",
          2871 => x"83",
          2872 => x"87",
          2873 => x"08",
          2874 => x"f1",
          2875 => x"c0",
          2876 => x"83",
          2877 => x"87",
          2878 => x"08",
          2879 => x"0c",
          2880 => x"8c",
          2881 => x"e0",
          2882 => x"83",
          2883 => x"80",
          2884 => x"9e",
          2885 => x"84",
          2886 => x"51",
          2887 => x"82",
          2888 => x"83",
          2889 => x"80",
          2890 => x"9e",
          2891 => x"88",
          2892 => x"51",
          2893 => x"80",
          2894 => x"81",
          2895 => x"f1",
          2896 => x"0b",
          2897 => x"90",
          2898 => x"80",
          2899 => x"52",
          2900 => x"2e",
          2901 => x"52",
          2902 => x"e7",
          2903 => x"87",
          2904 => x"08",
          2905 => x"80",
          2906 => x"52",
          2907 => x"83",
          2908 => x"71",
          2909 => x"34",
          2910 => x"c0",
          2911 => x"70",
          2912 => x"06",
          2913 => x"70",
          2914 => x"38",
          2915 => x"83",
          2916 => x"80",
          2917 => x"9e",
          2918 => x"90",
          2919 => x"51",
          2920 => x"80",
          2921 => x"81",
          2922 => x"f1",
          2923 => x"0b",
          2924 => x"90",
          2925 => x"80",
          2926 => x"52",
          2927 => x"2e",
          2928 => x"52",
          2929 => x"eb",
          2930 => x"87",
          2931 => x"08",
          2932 => x"80",
          2933 => x"52",
          2934 => x"83",
          2935 => x"71",
          2936 => x"34",
          2937 => x"c0",
          2938 => x"70",
          2939 => x"06",
          2940 => x"70",
          2941 => x"38",
          2942 => x"83",
          2943 => x"80",
          2944 => x"9e",
          2945 => x"80",
          2946 => x"51",
          2947 => x"80",
          2948 => x"81",
          2949 => x"f1",
          2950 => x"0b",
          2951 => x"90",
          2952 => x"80",
          2953 => x"52",
          2954 => x"83",
          2955 => x"71",
          2956 => x"34",
          2957 => x"90",
          2958 => x"06",
          2959 => x"53",
          2960 => x"f1",
          2961 => x"0b",
          2962 => x"90",
          2963 => x"80",
          2964 => x"52",
          2965 => x"83",
          2966 => x"71",
          2967 => x"34",
          2968 => x"90",
          2969 => x"06",
          2970 => x"53",
          2971 => x"f1",
          2972 => x"0b",
          2973 => x"90",
          2974 => x"06",
          2975 => x"70",
          2976 => x"38",
          2977 => x"83",
          2978 => x"87",
          2979 => x"08",
          2980 => x"70",
          2981 => x"34",
          2982 => x"04",
          2983 => x"82",
          2984 => x"0d",
          2985 => x"51",
          2986 => x"3f",
          2987 => x"33",
          2988 => x"aa",
          2989 => x"b4",
          2990 => x"3f",
          2991 => x"33",
          2992 => x"fa",
          2993 => x"eb",
          2994 => x"85",
          2995 => x"f1",
          2996 => x"75",
          2997 => x"83",
          2998 => x"55",
          2999 => x"38",
          3000 => x"33",
          3001 => x"d6",
          3002 => x"ef",
          3003 => x"84",
          3004 => x"f1",
          3005 => x"73",
          3006 => x"83",
          3007 => x"55",
          3008 => x"38",
          3009 => x"33",
          3010 => x"cf",
          3011 => x"e7",
          3012 => x"83",
          3013 => x"f1",
          3014 => x"74",
          3015 => x"83",
          3016 => x"56",
          3017 => x"38",
          3018 => x"33",
          3019 => x"ec",
          3020 => x"cc",
          3021 => x"3f",
          3022 => x"08",
          3023 => x"d8",
          3024 => x"c5",
          3025 => x"cc",
          3026 => x"d9",
          3027 => x"b5",
          3028 => x"f1",
          3029 => x"83",
          3030 => x"ff",
          3031 => x"83",
          3032 => x"c2",
          3033 => x"f1",
          3034 => x"83",
          3035 => x"ff",
          3036 => x"83",
          3037 => x"56",
          3038 => x"52",
          3039 => x"a6",
          3040 => x"e4",
          3041 => x"c0",
          3042 => x"31",
          3043 => x"b8",
          3044 => x"83",
          3045 => x"ff",
          3046 => x"83",
          3047 => x"55",
          3048 => x"38",
          3049 => x"33",
          3050 => x"38",
          3051 => x"af",
          3052 => x"0d",
          3053 => x"e0",
          3054 => x"84",
          3055 => x"51",
          3056 => x"84",
          3057 => x"bd",
          3058 => x"76",
          3059 => x"54",
          3060 => x"08",
          3061 => x"ac",
          3062 => x"ad",
          3063 => x"c2",
          3064 => x"3d",
          3065 => x"f1",
          3066 => x"bd",
          3067 => x"75",
          3068 => x"3f",
          3069 => x"08",
          3070 => x"29",
          3071 => x"54",
          3072 => x"e4",
          3073 => x"da",
          3074 => x"b3",
          3075 => x"f1",
          3076 => x"74",
          3077 => x"94",
          3078 => x"39",
          3079 => x"51",
          3080 => x"83",
          3081 => x"c0",
          3082 => x"f1",
          3083 => x"83",
          3084 => x"ff",
          3085 => x"83",
          3086 => x"52",
          3087 => x"51",
          3088 => x"3f",
          3089 => x"08",
          3090 => x"a8",
          3091 => x"b9",
          3092 => x"d0",
          3093 => x"3f",
          3094 => x"22",
          3095 => x"d8",
          3096 => x"a5",
          3097 => x"d8",
          3098 => x"84",
          3099 => x"51",
          3100 => x"84",
          3101 => x"bd",
          3102 => x"76",
          3103 => x"54",
          3104 => x"08",
          3105 => x"80",
          3106 => x"fd",
          3107 => x"eb",
          3108 => x"80",
          3109 => x"38",
          3110 => x"83",
          3111 => x"ff",
          3112 => x"83",
          3113 => x"54",
          3114 => x"fd",
          3115 => x"ec",
          3116 => x"94",
          3117 => x"bc",
          3118 => x"ed",
          3119 => x"80",
          3120 => x"38",
          3121 => x"db",
          3122 => x"bf",
          3123 => x"f1",
          3124 => x"74",
          3125 => x"c7",
          3126 => x"83",
          3127 => x"ff",
          3128 => x"83",
          3129 => x"54",
          3130 => x"fc",
          3131 => x"39",
          3132 => x"33",
          3133 => x"c0",
          3134 => x"8d",
          3135 => x"e5",
          3136 => x"80",
          3137 => x"38",
          3138 => x"f1",
          3139 => x"83",
          3140 => x"ff",
          3141 => x"83",
          3142 => x"55",
          3143 => x"fb",
          3144 => x"39",
          3145 => x"33",
          3146 => x"80",
          3147 => x"d9",
          3148 => x"f3",
          3149 => x"80",
          3150 => x"38",
          3151 => x"f1",
          3152 => x"f1",
          3153 => x"54",
          3154 => x"a0",
          3155 => x"b9",
          3156 => x"ef",
          3157 => x"80",
          3158 => x"38",
          3159 => x"f1",
          3160 => x"f1",
          3161 => x"54",
          3162 => x"bc",
          3163 => x"99",
          3164 => x"ea",
          3165 => x"80",
          3166 => x"38",
          3167 => x"f1",
          3168 => x"f1",
          3169 => x"54",
          3170 => x"d8",
          3171 => x"f9",
          3172 => x"e9",
          3173 => x"80",
          3174 => x"38",
          3175 => x"f1",
          3176 => x"f1",
          3177 => x"54",
          3178 => x"f4",
          3179 => x"d9",
          3180 => x"e8",
          3181 => x"80",
          3182 => x"38",
          3183 => x"f1",
          3184 => x"f1",
          3185 => x"54",
          3186 => x"90",
          3187 => x"b9",
          3188 => x"eb",
          3189 => x"80",
          3190 => x"38",
          3191 => x"dd",
          3192 => x"b0",
          3193 => x"d8",
          3194 => x"bd",
          3195 => x"f1",
          3196 => x"74",
          3197 => x"cd",
          3198 => x"ff",
          3199 => x"8e",
          3200 => x"71",
          3201 => x"38",
          3202 => x"83",
          3203 => x"52",
          3204 => x"83",
          3205 => x"ff",
          3206 => x"83",
          3207 => x"83",
          3208 => x"ff",
          3209 => x"83",
          3210 => x"83",
          3211 => x"ff",
          3212 => x"83",
          3213 => x"83",
          3214 => x"ff",
          3215 => x"83",
          3216 => x"83",
          3217 => x"ff",
          3218 => x"83",
          3219 => x"83",
          3220 => x"ff",
          3221 => x"83",
          3222 => x"71",
          3223 => x"04",
          3224 => x"c0",
          3225 => x"04",
          3226 => x"08",
          3227 => x"84",
          3228 => x"3d",
          3229 => x"08",
          3230 => x"5a",
          3231 => x"57",
          3232 => x"83",
          3233 => x"51",
          3234 => x"3f",
          3235 => x"08",
          3236 => x"8b",
          3237 => x"0b",
          3238 => x"08",
          3239 => x"f8",
          3240 => x"82",
          3241 => x"84",
          3242 => x"80",
          3243 => x"76",
          3244 => x"3f",
          3245 => x"08",
          3246 => x"55",
          3247 => x"b8",
          3248 => x"8e",
          3249 => x"e4",
          3250 => x"70",
          3251 => x"80",
          3252 => x"09",
          3253 => x"72",
          3254 => x"51",
          3255 => x"76",
          3256 => x"73",
          3257 => x"83",
          3258 => x"8c",
          3259 => x"51",
          3260 => x"3f",
          3261 => x"08",
          3262 => x"76",
          3263 => x"77",
          3264 => x"0c",
          3265 => x"04",
          3266 => x"51",
          3267 => x"3f",
          3268 => x"09",
          3269 => x"38",
          3270 => x"51",
          3271 => x"79",
          3272 => x"3f",
          3273 => x"56",
          3274 => x"08",
          3275 => x"52",
          3276 => x"51",
          3277 => x"3f",
          3278 => x"b8",
          3279 => x"3d",
          3280 => x"3d",
          3281 => x"08",
          3282 => x"71",
          3283 => x"33",
          3284 => x"57",
          3285 => x"81",
          3286 => x"0b",
          3287 => x"56",
          3288 => x"10",
          3289 => x"05",
          3290 => x"54",
          3291 => x"3f",
          3292 => x"08",
          3293 => x"73",
          3294 => x"9a",
          3295 => x"e4",
          3296 => x"84",
          3297 => x"73",
          3298 => x"88",
          3299 => x"2e",
          3300 => x"16",
          3301 => x"06",
          3302 => x"76",
          3303 => x"80",
          3304 => x"b8",
          3305 => x"3d",
          3306 => x"1a",
          3307 => x"ff",
          3308 => x"ff",
          3309 => x"c7",
          3310 => x"b8",
          3311 => x"2e",
          3312 => x"1b",
          3313 => x"76",
          3314 => x"3f",
          3315 => x"08",
          3316 => x"54",
          3317 => x"c9",
          3318 => x"70",
          3319 => x"57",
          3320 => x"27",
          3321 => x"ff",
          3322 => x"33",
          3323 => x"76",
          3324 => x"e6",
          3325 => x"70",
          3326 => x"55",
          3327 => x"2e",
          3328 => x"fe",
          3329 => x"75",
          3330 => x"80",
          3331 => x"59",
          3332 => x"39",
          3333 => x"e4",
          3334 => x"f2",
          3335 => x"56",
          3336 => x"3f",
          3337 => x"08",
          3338 => x"83",
          3339 => x"53",
          3340 => x"77",
          3341 => x"fd",
          3342 => x"e4",
          3343 => x"ba",
          3344 => x"ff",
          3345 => x"84",
          3346 => x"55",
          3347 => x"b8",
          3348 => x"9d",
          3349 => x"e4",
          3350 => x"70",
          3351 => x"80",
          3352 => x"53",
          3353 => x"16",
          3354 => x"52",
          3355 => x"99",
          3356 => x"2e",
          3357 => x"ff",
          3358 => x"0b",
          3359 => x"0c",
          3360 => x"04",
          3361 => x"b5",
          3362 => x"3d",
          3363 => x"08",
          3364 => x"80",
          3365 => x"34",
          3366 => x"33",
          3367 => x"08",
          3368 => x"9e",
          3369 => x"f2",
          3370 => x"56",
          3371 => x"82",
          3372 => x"80",
          3373 => x"38",
          3374 => x"06",
          3375 => x"90",
          3376 => x"80",
          3377 => x"38",
          3378 => x"3d",
          3379 => x"51",
          3380 => x"84",
          3381 => x"98",
          3382 => x"2c",
          3383 => x"ff",
          3384 => x"79",
          3385 => x"84",
          3386 => x"70",
          3387 => x"98",
          3388 => x"9c",
          3389 => x"2b",
          3390 => x"71",
          3391 => x"70",
          3392 => x"dd",
          3393 => x"08",
          3394 => x"52",
          3395 => x"46",
          3396 => x"5c",
          3397 => x"74",
          3398 => x"cd",
          3399 => x"27",
          3400 => x"75",
          3401 => x"29",
          3402 => x"05",
          3403 => x"57",
          3404 => x"24",
          3405 => x"75",
          3406 => x"82",
          3407 => x"80",
          3408 => x"f0",
          3409 => x"57",
          3410 => x"91",
          3411 => x"ec",
          3412 => x"70",
          3413 => x"78",
          3414 => x"95",
          3415 => x"2e",
          3416 => x"84",
          3417 => x"81",
          3418 => x"2e",
          3419 => x"81",
          3420 => x"2b",
          3421 => x"84",
          3422 => x"70",
          3423 => x"97",
          3424 => x"2c",
          3425 => x"2b",
          3426 => x"11",
          3427 => x"5f",
          3428 => x"57",
          3429 => x"2e",
          3430 => x"76",
          3431 => x"34",
          3432 => x"81",
          3433 => x"ba",
          3434 => x"80",
          3435 => x"80",
          3436 => x"98",
          3437 => x"ff",
          3438 => x"41",
          3439 => x"80",
          3440 => x"10",
          3441 => x"2b",
          3442 => x"0b",
          3443 => x"16",
          3444 => x"77",
          3445 => x"38",
          3446 => x"15",
          3447 => x"33",
          3448 => x"61",
          3449 => x"38",
          3450 => x"ff",
          3451 => x"f2",
          3452 => x"76",
          3453 => x"ab",
          3454 => x"39",
          3455 => x"b2",
          3456 => x"76",
          3457 => x"76",
          3458 => x"34",
          3459 => x"9c",
          3460 => x"34",
          3461 => x"62",
          3462 => x"26",
          3463 => x"74",
          3464 => x"c3",
          3465 => x"76",
          3466 => x"dd",
          3467 => x"7f",
          3468 => x"84",
          3469 => x"80",
          3470 => x"9c",
          3471 => x"84",
          3472 => x"56",
          3473 => x"fd",
          3474 => x"d4",
          3475 => x"88",
          3476 => x"9b",
          3477 => x"a8",
          3478 => x"57",
          3479 => x"a8",
          3480 => x"39",
          3481 => x"33",
          3482 => x"06",
          3483 => x"33",
          3484 => x"75",
          3485 => x"d6",
          3486 => x"c8",
          3487 => x"15",
          3488 => x"d0",
          3489 => x"16",
          3490 => x"55",
          3491 => x"3f",
          3492 => x"7c",
          3493 => x"da",
          3494 => x"10",
          3495 => x"05",
          3496 => x"59",
          3497 => x"38",
          3498 => x"a4",
          3499 => x"34",
          3500 => x"33",
          3501 => x"33",
          3502 => x"80",
          3503 => x"84",
          3504 => x"52",
          3505 => x"b5",
          3506 => x"d4",
          3507 => x"a0",
          3508 => x"9b",
          3509 => x"c8",
          3510 => x"51",
          3511 => x"3f",
          3512 => x"33",
          3513 => x"7a",
          3514 => x"34",
          3515 => x"06",
          3516 => x"38",
          3517 => x"a6",
          3518 => x"84",
          3519 => x"fb",
          3520 => x"8a",
          3521 => x"c8",
          3522 => x"8d",
          3523 => x"10",
          3524 => x"fc",
          3525 => x"08",
          3526 => x"8e",
          3527 => x"08",
          3528 => x"2e",
          3529 => x"75",
          3530 => x"fd",
          3531 => x"e4",
          3532 => x"a4",
          3533 => x"e4",
          3534 => x"06",
          3535 => x"75",
          3536 => x"ff",
          3537 => x"84",
          3538 => x"84",
          3539 => x"56",
          3540 => x"2e",
          3541 => x"84",
          3542 => x"52",
          3543 => x"b4",
          3544 => x"d4",
          3545 => x"a0",
          3546 => x"83",
          3547 => x"c8",
          3548 => x"51",
          3549 => x"3f",
          3550 => x"33",
          3551 => x"74",
          3552 => x"34",
          3553 => x"06",
          3554 => x"84",
          3555 => x"70",
          3556 => x"84",
          3557 => x"5b",
          3558 => x"79",
          3559 => x"38",
          3560 => x"08",
          3561 => x"57",
          3562 => x"a8",
          3563 => x"70",
          3564 => x"ff",
          3565 => x"84",
          3566 => x"70",
          3567 => x"84",
          3568 => x"5a",
          3569 => x"78",
          3570 => x"38",
          3571 => x"08",
          3572 => x"57",
          3573 => x"a8",
          3574 => x"70",
          3575 => x"ff",
          3576 => x"84",
          3577 => x"70",
          3578 => x"84",
          3579 => x"5a",
          3580 => x"76",
          3581 => x"38",
          3582 => x"84",
          3583 => x"84",
          3584 => x"56",
          3585 => x"2e",
          3586 => x"ff",
          3587 => x"84",
          3588 => x"75",
          3589 => x"98",
          3590 => x"ff",
          3591 => x"5a",
          3592 => x"80",
          3593 => x"d4",
          3594 => x"a0",
          3595 => x"bf",
          3596 => x"a8",
          3597 => x"2b",
          3598 => x"84",
          3599 => x"5a",
          3600 => x"74",
          3601 => x"86",
          3602 => x"c8",
          3603 => x"51",
          3604 => x"3f",
          3605 => x"0a",
          3606 => x"0a",
          3607 => x"2c",
          3608 => x"33",
          3609 => x"74",
          3610 => x"e2",
          3611 => x"c8",
          3612 => x"51",
          3613 => x"3f",
          3614 => x"0a",
          3615 => x"0a",
          3616 => x"2c",
          3617 => x"33",
          3618 => x"7a",
          3619 => x"b9",
          3620 => x"39",
          3621 => x"81",
          3622 => x"34",
          3623 => x"08",
          3624 => x"51",
          3625 => x"3f",
          3626 => x"0a",
          3627 => x"0a",
          3628 => x"2c",
          3629 => x"33",
          3630 => x"75",
          3631 => x"e6",
          3632 => x"58",
          3633 => x"78",
          3634 => x"c8",
          3635 => x"33",
          3636 => x"9b",
          3637 => x"80",
          3638 => x"80",
          3639 => x"98",
          3640 => x"a4",
          3641 => x"55",
          3642 => x"ff",
          3643 => x"b6",
          3644 => x"a8",
          3645 => x"80",
          3646 => x"38",
          3647 => x"08",
          3648 => x"ff",
          3649 => x"84",
          3650 => x"ff",
          3651 => x"84",
          3652 => x"76",
          3653 => x"55",
          3654 => x"d0",
          3655 => x"05",
          3656 => x"34",
          3657 => x"08",
          3658 => x"ff",
          3659 => x"84",
          3660 => x"7b",
          3661 => x"3f",
          3662 => x"08",
          3663 => x"58",
          3664 => x"38",
          3665 => x"33",
          3666 => x"2e",
          3667 => x"83",
          3668 => x"70",
          3669 => x"f1",
          3670 => x"08",
          3671 => x"74",
          3672 => x"75",
          3673 => x"fc",
          3674 => x"fc",
          3675 => x"70",
          3676 => x"80",
          3677 => x"84",
          3678 => x"7b",
          3679 => x"d4",
          3680 => x"10",
          3681 => x"05",
          3682 => x"41",
          3683 => x"ad",
          3684 => x"d0",
          3685 => x"80",
          3686 => x"83",
          3687 => x"58",
          3688 => x"8b",
          3689 => x"0b",
          3690 => x"34",
          3691 => x"d0",
          3692 => x"84",
          3693 => x"b4",
          3694 => x"84",
          3695 => x"55",
          3696 => x"b6",
          3697 => x"c8",
          3698 => x"51",
          3699 => x"3f",
          3700 => x"08",
          3701 => x"ff",
          3702 => x"84",
          3703 => x"52",
          3704 => x"af",
          3705 => x"d0",
          3706 => x"05",
          3707 => x"d0",
          3708 => x"81",
          3709 => x"74",
          3710 => x"d1",
          3711 => x"a0",
          3712 => x"0b",
          3713 => x"34",
          3714 => x"d0",
          3715 => x"be",
          3716 => x"34",
          3717 => x"1d",
          3718 => x"a8",
          3719 => x"80",
          3720 => x"84",
          3721 => x"52",
          3722 => x"ae",
          3723 => x"d4",
          3724 => x"a0",
          3725 => x"b7",
          3726 => x"c8",
          3727 => x"51",
          3728 => x"3f",
          3729 => x"33",
          3730 => x"7c",
          3731 => x"34",
          3732 => x"06",
          3733 => x"38",
          3734 => x"51",
          3735 => x"3f",
          3736 => x"d0",
          3737 => x"0b",
          3738 => x"34",
          3739 => x"e4",
          3740 => x"0d",
          3741 => x"a8",
          3742 => x"ff",
          3743 => x"7a",
          3744 => x"ca",
          3745 => x"a4",
          3746 => x"59",
          3747 => x"a4",
          3748 => x"58",
          3749 => x"a8",
          3750 => x"c8",
          3751 => x"51",
          3752 => x"3f",
          3753 => x"33",
          3754 => x"70",
          3755 => x"d0",
          3756 => x"52",
          3757 => x"76",
          3758 => x"38",
          3759 => x"08",
          3760 => x"ff",
          3761 => x"84",
          3762 => x"70",
          3763 => x"98",
          3764 => x"a4",
          3765 => x"59",
          3766 => x"24",
          3767 => x"84",
          3768 => x"52",
          3769 => x"ad",
          3770 => x"81",
          3771 => x"81",
          3772 => x"70",
          3773 => x"d0",
          3774 => x"51",
          3775 => x"24",
          3776 => x"84",
          3777 => x"52",
          3778 => x"ac",
          3779 => x"81",
          3780 => x"81",
          3781 => x"70",
          3782 => x"d0",
          3783 => x"51",
          3784 => x"25",
          3785 => x"f3",
          3786 => x"16",
          3787 => x"33",
          3788 => x"d4",
          3789 => x"76",
          3790 => x"ac",
          3791 => x"81",
          3792 => x"81",
          3793 => x"70",
          3794 => x"d0",
          3795 => x"57",
          3796 => x"25",
          3797 => x"7b",
          3798 => x"17",
          3799 => x"84",
          3800 => x"52",
          3801 => x"ff",
          3802 => x"75",
          3803 => x"29",
          3804 => x"05",
          3805 => x"84",
          3806 => x"43",
          3807 => x"76",
          3808 => x"38",
          3809 => x"84",
          3810 => x"70",
          3811 => x"58",
          3812 => x"2e",
          3813 => x"84",
          3814 => x"55",
          3815 => x"ae",
          3816 => x"2b",
          3817 => x"57",
          3818 => x"24",
          3819 => x"16",
          3820 => x"81",
          3821 => x"81",
          3822 => x"81",
          3823 => x"70",
          3824 => x"d0",
          3825 => x"57",
          3826 => x"25",
          3827 => x"18",
          3828 => x"d0",
          3829 => x"81",
          3830 => x"05",
          3831 => x"33",
          3832 => x"d0",
          3833 => x"76",
          3834 => x"38",
          3835 => x"75",
          3836 => x"34",
          3837 => x"d0",
          3838 => x"81",
          3839 => x"81",
          3840 => x"70",
          3841 => x"81",
          3842 => x"58",
          3843 => x"76",
          3844 => x"38",
          3845 => x"70",
          3846 => x"81",
          3847 => x"57",
          3848 => x"25",
          3849 => x"84",
          3850 => x"52",
          3851 => x"aa",
          3852 => x"81",
          3853 => x"81",
          3854 => x"70",
          3855 => x"d0",
          3856 => x"57",
          3857 => x"25",
          3858 => x"84",
          3859 => x"52",
          3860 => x"aa",
          3861 => x"81",
          3862 => x"81",
          3863 => x"70",
          3864 => x"d0",
          3865 => x"57",
          3866 => x"24",
          3867 => x"f0",
          3868 => x"f1",
          3869 => x"75",
          3870 => x"9d",
          3871 => x"ff",
          3872 => x"84",
          3873 => x"84",
          3874 => x"84",
          3875 => x"81",
          3876 => x"05",
          3877 => x"7b",
          3878 => x"cf",
          3879 => x"a4",
          3880 => x"a8",
          3881 => x"74",
          3882 => x"c8",
          3883 => x"c8",
          3884 => x"51",
          3885 => x"3f",
          3886 => x"08",
          3887 => x"ff",
          3888 => x"84",
          3889 => x"52",
          3890 => x"a9",
          3891 => x"d0",
          3892 => x"05",
          3893 => x"d0",
          3894 => x"81",
          3895 => x"c7",
          3896 => x"80",
          3897 => x"84",
          3898 => x"83",
          3899 => x"84",
          3900 => x"85",
          3901 => x"83",
          3902 => x"77",
          3903 => x"80",
          3904 => x"d4",
          3905 => x"7b",
          3906 => x"52",
          3907 => x"df",
          3908 => x"80",
          3909 => x"80",
          3910 => x"98",
          3911 => x"a4",
          3912 => x"57",
          3913 => x"da",
          3914 => x"a8",
          3915 => x"2b",
          3916 => x"79",
          3917 => x"5d",
          3918 => x"75",
          3919 => x"8e",
          3920 => x"39",
          3921 => x"08",
          3922 => x"fc",
          3923 => x"fc",
          3924 => x"76",
          3925 => x"bb",
          3926 => x"84",
          3927 => x"75",
          3928 => x"38",
          3929 => x"f2",
          3930 => x"f2",
          3931 => x"74",
          3932 => x"d4",
          3933 => x"81",
          3934 => x"83",
          3935 => x"51",
          3936 => x"3f",
          3937 => x"f2",
          3938 => x"3d",
          3939 => x"5f",
          3940 => x"74",
          3941 => x"e9",
          3942 => x"0c",
          3943 => x"18",
          3944 => x"80",
          3945 => x"38",
          3946 => x"75",
          3947 => x"f9",
          3948 => x"e4",
          3949 => x"a4",
          3950 => x"e4",
          3951 => x"06",
          3952 => x"75",
          3953 => x"ff",
          3954 => x"93",
          3955 => x"a4",
          3956 => x"a8",
          3957 => x"5d",
          3958 => x"f2",
          3959 => x"d4",
          3960 => x"88",
          3961 => x"87",
          3962 => x"c8",
          3963 => x"51",
          3964 => x"3f",
          3965 => x"08",
          3966 => x"ff",
          3967 => x"84",
          3968 => x"ff",
          3969 => x"84",
          3970 => x"79",
          3971 => x"55",
          3972 => x"7c",
          3973 => x"84",
          3974 => x"80",
          3975 => x"a4",
          3976 => x"b8",
          3977 => x"3d",
          3978 => x"51",
          3979 => x"3f",
          3980 => x"08",
          3981 => x"34",
          3982 => x"08",
          3983 => x"81",
          3984 => x"52",
          3985 => x"aa",
          3986 => x"1d",
          3987 => x"06",
          3988 => x"33",
          3989 => x"33",
          3990 => x"56",
          3991 => x"f1",
          3992 => x"d4",
          3993 => x"88",
          3994 => x"83",
          3995 => x"c8",
          3996 => x"51",
          3997 => x"3f",
          3998 => x"08",
          3999 => x"ff",
          4000 => x"84",
          4001 => x"ff",
          4002 => x"84",
          4003 => x"76",
          4004 => x"55",
          4005 => x"51",
          4006 => x"3f",
          4007 => x"08",
          4008 => x"34",
          4009 => x"08",
          4010 => x"81",
          4011 => x"52",
          4012 => x"a9",
          4013 => x"1d",
          4014 => x"06",
          4015 => x"33",
          4016 => x"33",
          4017 => x"58",
          4018 => x"f0",
          4019 => x"d4",
          4020 => x"88",
          4021 => x"97",
          4022 => x"c8",
          4023 => x"51",
          4024 => x"3f",
          4025 => x"08",
          4026 => x"ff",
          4027 => x"84",
          4028 => x"ff",
          4029 => x"84",
          4030 => x"60",
          4031 => x"55",
          4032 => x"51",
          4033 => x"3f",
          4034 => x"33",
          4035 => x"87",
          4036 => x"f1",
          4037 => x"19",
          4038 => x"5c",
          4039 => x"d1",
          4040 => x"e4",
          4041 => x"83",
          4042 => x"70",
          4043 => x"f1",
          4044 => x"08",
          4045 => x"74",
          4046 => x"d5",
          4047 => x"7b",
          4048 => x"ff",
          4049 => x"83",
          4050 => x"81",
          4051 => x"ff",
          4052 => x"93",
          4053 => x"f2",
          4054 => x"f2",
          4055 => x"b1",
          4056 => x"fe",
          4057 => x"76",
          4058 => x"75",
          4059 => x"c0",
          4060 => x"d0",
          4061 => x"51",
          4062 => x"3f",
          4063 => x"08",
          4064 => x"f3",
          4065 => x"84",
          4066 => x"80",
          4067 => x"a4",
          4068 => x"b8",
          4069 => x"3d",
          4070 => x"53",
          4071 => x"b8",
          4072 => x"81",
          4073 => x"84",
          4074 => x"82",
          4075 => x"b8",
          4076 => x"3d",
          4077 => x"f2",
          4078 => x"80",
          4079 => x"51",
          4080 => x"3f",
          4081 => x"08",
          4082 => x"e4",
          4083 => x"09",
          4084 => x"ee",
          4085 => x"e4",
          4086 => x"a6",
          4087 => x"b8",
          4088 => x"80",
          4089 => x"e4",
          4090 => x"e3",
          4091 => x"e4",
          4092 => x"70",
          4093 => x"80",
          4094 => x"81",
          4095 => x"f2",
          4096 => x"10",
          4097 => x"fc",
          4098 => x"58",
          4099 => x"74",
          4100 => x"76",
          4101 => x"fc",
          4102 => x"fc",
          4103 => x"70",
          4104 => x"80",
          4105 => x"84",
          4106 => x"75",
          4107 => x"d4",
          4108 => x"10",
          4109 => x"05",
          4110 => x"40",
          4111 => x"38",
          4112 => x"81",
          4113 => x"57",
          4114 => x"83",
          4115 => x"75",
          4116 => x"81",
          4117 => x"38",
          4118 => x"38",
          4119 => x"76",
          4120 => x"74",
          4121 => x"83",
          4122 => x"d4",
          4123 => x"70",
          4124 => x"5b",
          4125 => x"27",
          4126 => x"80",
          4127 => x"d4",
          4128 => x"39",
          4129 => x"d3",
          4130 => x"f2",
          4131 => x"82",
          4132 => x"06",
          4133 => x"05",
          4134 => x"54",
          4135 => x"80",
          4136 => x"84",
          4137 => x"75",
          4138 => x"d4",
          4139 => x"10",
          4140 => x"05",
          4141 => x"40",
          4142 => x"2e",
          4143 => x"ff",
          4144 => x"83",
          4145 => x"fe",
          4146 => x"83",
          4147 => x"f1",
          4148 => x"e0",
          4149 => x"9f",
          4150 => x"e7",
          4151 => x"e4",
          4152 => x"0d",
          4153 => x"05",
          4154 => x"05",
          4155 => x"33",
          4156 => x"83",
          4157 => x"38",
          4158 => x"81",
          4159 => x"73",
          4160 => x"38",
          4161 => x"82",
          4162 => x"a7",
          4163 => x"86",
          4164 => x"70",
          4165 => x"56",
          4166 => x"79",
          4167 => x"38",
          4168 => x"94",
          4169 => x"f8",
          4170 => x"83",
          4171 => x"83",
          4172 => x"70",
          4173 => x"90",
          4174 => x"88",
          4175 => x"07",
          4176 => x"56",
          4177 => x"77",
          4178 => x"80",
          4179 => x"05",
          4180 => x"73",
          4181 => x"55",
          4182 => x"26",
          4183 => x"78",
          4184 => x"83",
          4185 => x"84",
          4186 => x"79",
          4187 => x"55",
          4188 => x"e0",
          4189 => x"74",
          4190 => x"05",
          4191 => x"13",
          4192 => x"38",
          4193 => x"04",
          4194 => x"80",
          4195 => x"94",
          4196 => x"10",
          4197 => x"95",
          4198 => x"29",
          4199 => x"5b",
          4200 => x"59",
          4201 => x"80",
          4202 => x"d8",
          4203 => x"ff",
          4204 => x"d7",
          4205 => x"ff",
          4206 => x"92",
          4207 => x"ff",
          4208 => x"75",
          4209 => x"5d",
          4210 => x"5b",
          4211 => x"26",
          4212 => x"74",
          4213 => x"56",
          4214 => x"06",
          4215 => x"06",
          4216 => x"06",
          4217 => x"ff",
          4218 => x"ff",
          4219 => x"29",
          4220 => x"57",
          4221 => x"74",
          4222 => x"38",
          4223 => x"33",
          4224 => x"05",
          4225 => x"1b",
          4226 => x"83",
          4227 => x"80",
          4228 => x"38",
          4229 => x"53",
          4230 => x"fe",
          4231 => x"73",
          4232 => x"55",
          4233 => x"90",
          4234 => x"81",
          4235 => x"e8",
          4236 => x"a0",
          4237 => x"a7",
          4238 => x"84",
          4239 => x"70",
          4240 => x"84",
          4241 => x"70",
          4242 => x"83",
          4243 => x"70",
          4244 => x"5b",
          4245 => x"56",
          4246 => x"78",
          4247 => x"38",
          4248 => x"06",
          4249 => x"06",
          4250 => x"18",
          4251 => x"79",
          4252 => x"bb",
          4253 => x"83",
          4254 => x"80",
          4255 => x"95",
          4256 => x"90",
          4257 => x"2b",
          4258 => x"07",
          4259 => x"07",
          4260 => x"7f",
          4261 => x"5b",
          4262 => x"fd",
          4263 => x"be",
          4264 => x"e6",
          4265 => x"94",
          4266 => x"ff",
          4267 => x"10",
          4268 => x"95",
          4269 => x"29",
          4270 => x"a0",
          4271 => x"57",
          4272 => x"5f",
          4273 => x"80",
          4274 => x"b6",
          4275 => x"81",
          4276 => x"b6",
          4277 => x"81",
          4278 => x"f8",
          4279 => x"83",
          4280 => x"7c",
          4281 => x"05",
          4282 => x"5f",
          4283 => x"5e",
          4284 => x"26",
          4285 => x"7a",
          4286 => x"7d",
          4287 => x"53",
          4288 => x"06",
          4289 => x"06",
          4290 => x"7d",
          4291 => x"06",
          4292 => x"06",
          4293 => x"58",
          4294 => x"5d",
          4295 => x"26",
          4296 => x"75",
          4297 => x"73",
          4298 => x"83",
          4299 => x"79",
          4300 => x"76",
          4301 => x"7b",
          4302 => x"fb",
          4303 => x"78",
          4304 => x"56",
          4305 => x"fb",
          4306 => x"ee",
          4307 => x"ff",
          4308 => x"87",
          4309 => x"73",
          4310 => x"34",
          4311 => x"9c",
          4312 => x"75",
          4313 => x"75",
          4314 => x"80",
          4315 => x"76",
          4316 => x"34",
          4317 => x"94",
          4318 => x"34",
          4319 => x"ff",
          4320 => x"81",
          4321 => x"fa",
          4322 => x"a0",
          4323 => x"08",
          4324 => x"f8",
          4325 => x"81",
          4326 => x"06",
          4327 => x"55",
          4328 => x"73",
          4329 => x"ff",
          4330 => x"07",
          4331 => x"75",
          4332 => x"87",
          4333 => x"77",
          4334 => x"51",
          4335 => x"a0",
          4336 => x"73",
          4337 => x"06",
          4338 => x"72",
          4339 => x"d0",
          4340 => x"d8",
          4341 => x"84",
          4342 => x"87",
          4343 => x"84",
          4344 => x"84",
          4345 => x"04",
          4346 => x"02",
          4347 => x"02",
          4348 => x"05",
          4349 => x"d7",
          4350 => x"56",
          4351 => x"79",
          4352 => x"38",
          4353 => x"33",
          4354 => x"33",
          4355 => x"33",
          4356 => x"12",
          4357 => x"80",
          4358 => x"92",
          4359 => x"57",
          4360 => x"29",
          4361 => x"ff",
          4362 => x"f6",
          4363 => x"57",
          4364 => x"81",
          4365 => x"38",
          4366 => x"22",
          4367 => x"74",
          4368 => x"23",
          4369 => x"33",
          4370 => x"81",
          4371 => x"81",
          4372 => x"5b",
          4373 => x"26",
          4374 => x"ff",
          4375 => x"83",
          4376 => x"83",
          4377 => x"70",
          4378 => x"06",
          4379 => x"33",
          4380 => x"79",
          4381 => x"89",
          4382 => x"d8",
          4383 => x"29",
          4384 => x"54",
          4385 => x"26",
          4386 => x"97",
          4387 => x"54",
          4388 => x"13",
          4389 => x"16",
          4390 => x"81",
          4391 => x"75",
          4392 => x"57",
          4393 => x"54",
          4394 => x"73",
          4395 => x"73",
          4396 => x"a1",
          4397 => x"90",
          4398 => x"b6",
          4399 => x"a0",
          4400 => x"14",
          4401 => x"70",
          4402 => x"34",
          4403 => x"9f",
          4404 => x"eb",
          4405 => x"d6",
          4406 => x"56",
          4407 => x"92",
          4408 => x"78",
          4409 => x"77",
          4410 => x"06",
          4411 => x"73",
          4412 => x"38",
          4413 => x"81",
          4414 => x"d8",
          4415 => x"29",
          4416 => x"75",
          4417 => x"a0",
          4418 => x"a7",
          4419 => x"81",
          4420 => x"81",
          4421 => x"71",
          4422 => x"5c",
          4423 => x"79",
          4424 => x"84",
          4425 => x"54",
          4426 => x"33",
          4427 => x"e0",
          4428 => x"70",
          4429 => x"34",
          4430 => x"05",
          4431 => x"70",
          4432 => x"34",
          4433 => x"b6",
          4434 => x"b6",
          4435 => x"71",
          4436 => x"5c",
          4437 => x"75",
          4438 => x"80",
          4439 => x"b8",
          4440 => x"3d",
          4441 => x"83",
          4442 => x"83",
          4443 => x"70",
          4444 => x"06",
          4445 => x"33",
          4446 => x"73",
          4447 => x"f9",
          4448 => x"2e",
          4449 => x"78",
          4450 => x"ff",
          4451 => x"94",
          4452 => x"72",
          4453 => x"81",
          4454 => x"38",
          4455 => x"81",
          4456 => x"d8",
          4457 => x"29",
          4458 => x"11",
          4459 => x"54",
          4460 => x"fe",
          4461 => x"f8",
          4462 => x"97",
          4463 => x"76",
          4464 => x"56",
          4465 => x"e0",
          4466 => x"75",
          4467 => x"57",
          4468 => x"53",
          4469 => x"fe",
          4470 => x"0b",
          4471 => x"34",
          4472 => x"81",
          4473 => x"ff",
          4474 => x"d8",
          4475 => x"39",
          4476 => x"b6",
          4477 => x"56",
          4478 => x"83",
          4479 => x"33",
          4480 => x"e0",
          4481 => x"34",
          4482 => x"33",
          4483 => x"39",
          4484 => x"76",
          4485 => x"9f",
          4486 => x"51",
          4487 => x"9b",
          4488 => x"10",
          4489 => x"05",
          4490 => x"04",
          4491 => x"33",
          4492 => x"27",
          4493 => x"83",
          4494 => x"80",
          4495 => x"e4",
          4496 => x"0d",
          4497 => x"83",
          4498 => x"83",
          4499 => x"70",
          4500 => x"54",
          4501 => x"2e",
          4502 => x"12",
          4503 => x"f8",
          4504 => x"0b",
          4505 => x"0c",
          4506 => x"04",
          4507 => x"33",
          4508 => x"70",
          4509 => x"2c",
          4510 => x"55",
          4511 => x"83",
          4512 => x"de",
          4513 => x"94",
          4514 => x"84",
          4515 => x"ff",
          4516 => x"51",
          4517 => x"83",
          4518 => x"72",
          4519 => x"34",
          4520 => x"b8",
          4521 => x"3d",
          4522 => x"f8",
          4523 => x"73",
          4524 => x"70",
          4525 => x"06",
          4526 => x"55",
          4527 => x"95",
          4528 => x"84",
          4529 => x"86",
          4530 => x"83",
          4531 => x"72",
          4532 => x"d8",
          4533 => x"55",
          4534 => x"74",
          4535 => x"70",
          4536 => x"f8",
          4537 => x"0b",
          4538 => x"0c",
          4539 => x"04",
          4540 => x"f8",
          4541 => x"f8",
          4542 => x"b6",
          4543 => x"05",
          4544 => x"75",
          4545 => x"38",
          4546 => x"70",
          4547 => x"34",
          4548 => x"ff",
          4549 => x"8f",
          4550 => x"70",
          4551 => x"38",
          4552 => x"83",
          4553 => x"51",
          4554 => x"83",
          4555 => x"70",
          4556 => x"71",
          4557 => x"f0",
          4558 => x"84",
          4559 => x"52",
          4560 => x"80",
          4561 => x"81",
          4562 => x"80",
          4563 => x"f8",
          4564 => x"0b",
          4565 => x"0c",
          4566 => x"04",
          4567 => x"33",
          4568 => x"90",
          4569 => x"83",
          4570 => x"80",
          4571 => x"e4",
          4572 => x"0d",
          4573 => x"90",
          4574 => x"07",
          4575 => x"f8",
          4576 => x"39",
          4577 => x"33",
          4578 => x"86",
          4579 => x"83",
          4580 => x"d7",
          4581 => x"0b",
          4582 => x"34",
          4583 => x"b8",
          4584 => x"3d",
          4585 => x"f8",
          4586 => x"fc",
          4587 => x"51",
          4588 => x"90",
          4589 => x"39",
          4590 => x"33",
          4591 => x"70",
          4592 => x"34",
          4593 => x"83",
          4594 => x"81",
          4595 => x"07",
          4596 => x"f8",
          4597 => x"93",
          4598 => x"90",
          4599 => x"06",
          4600 => x"70",
          4601 => x"34",
          4602 => x"83",
          4603 => x"81",
          4604 => x"07",
          4605 => x"f8",
          4606 => x"ef",
          4607 => x"90",
          4608 => x"06",
          4609 => x"f8",
          4610 => x"df",
          4611 => x"90",
          4612 => x"06",
          4613 => x"51",
          4614 => x"90",
          4615 => x"39",
          4616 => x"33",
          4617 => x"b0",
          4618 => x"83",
          4619 => x"fe",
          4620 => x"f8",
          4621 => x"ef",
          4622 => x"07",
          4623 => x"f8",
          4624 => x"a7",
          4625 => x"90",
          4626 => x"06",
          4627 => x"51",
          4628 => x"90",
          4629 => x"39",
          4630 => x"33",
          4631 => x"a0",
          4632 => x"83",
          4633 => x"fe",
          4634 => x"f8",
          4635 => x"8f",
          4636 => x"83",
          4637 => x"fd",
          4638 => x"f8",
          4639 => x"fa",
          4640 => x"51",
          4641 => x"90",
          4642 => x"39",
          4643 => x"02",
          4644 => x"02",
          4645 => x"c3",
          4646 => x"f8",
          4647 => x"f8",
          4648 => x"f8",
          4649 => x"b6",
          4650 => x"41",
          4651 => x"59",
          4652 => x"82",
          4653 => x"82",
          4654 => x"78",
          4655 => x"82",
          4656 => x"b6",
          4657 => x"0b",
          4658 => x"34",
          4659 => x"94",
          4660 => x"f8",
          4661 => x"83",
          4662 => x"8f",
          4663 => x"78",
          4664 => x"81",
          4665 => x"80",
          4666 => x"da",
          4667 => x"84",
          4668 => x"82",
          4669 => x"94",
          4670 => x"83",
          4671 => x"82",
          4672 => x"92",
          4673 => x"84",
          4674 => x"57",
          4675 => x"33",
          4676 => x"d6",
          4677 => x"54",
          4678 => x"52",
          4679 => x"51",
          4680 => x"3f",
          4681 => x"da",
          4682 => x"84",
          4683 => x"7a",
          4684 => x"34",
          4685 => x"92",
          4686 => x"f8",
          4687 => x"3d",
          4688 => x"0b",
          4689 => x"34",
          4690 => x"b6",
          4691 => x"0b",
          4692 => x"34",
          4693 => x"f8",
          4694 => x"0b",
          4695 => x"23",
          4696 => x"33",
          4697 => x"e6",
          4698 => x"b7",
          4699 => x"79",
          4700 => x"7c",
          4701 => x"83",
          4702 => x"ff",
          4703 => x"80",
          4704 => x"e5",
          4705 => x"79",
          4706 => x"38",
          4707 => x"b8",
          4708 => x"22",
          4709 => x"e3",
          4710 => x"80",
          4711 => x"1a",
          4712 => x"06",
          4713 => x"33",
          4714 => x"78",
          4715 => x"38",
          4716 => x"51",
          4717 => x"3f",
          4718 => x"da",
          4719 => x"84",
          4720 => x"7a",
          4721 => x"34",
          4722 => x"92",
          4723 => x"f8",
          4724 => x"3d",
          4725 => x"0b",
          4726 => x"34",
          4727 => x"b6",
          4728 => x"0b",
          4729 => x"34",
          4730 => x"f8",
          4731 => x"0b",
          4732 => x"23",
          4733 => x"51",
          4734 => x"3f",
          4735 => x"08",
          4736 => x"90",
          4737 => x"81",
          4738 => x"83",
          4739 => x"ff",
          4740 => x"78",
          4741 => x"08",
          4742 => x"38",
          4743 => x"19",
          4744 => x"e3",
          4745 => x"ff",
          4746 => x"19",
          4747 => x"06",
          4748 => x"39",
          4749 => x"7a",
          4750 => x"a7",
          4751 => x"b6",
          4752 => x"f8",
          4753 => x"f8",
          4754 => x"71",
          4755 => x"a7",
          4756 => x"83",
          4757 => x"53",
          4758 => x"71",
          4759 => x"70",
          4760 => x"06",
          4761 => x"33",
          4762 => x"55",
          4763 => x"81",
          4764 => x"38",
          4765 => x"81",
          4766 => x"89",
          4767 => x"38",
          4768 => x"83",
          4769 => x"88",
          4770 => x"38",
          4771 => x"33",
          4772 => x"33",
          4773 => x"33",
          4774 => x"05",
          4775 => x"84",
          4776 => x"33",
          4777 => x"80",
          4778 => x"b6",
          4779 => x"f8",
          4780 => x"f8",
          4781 => x"71",
          4782 => x"5a",
          4783 => x"83",
          4784 => x"34",
          4785 => x"33",
          4786 => x"16",
          4787 => x"f8",
          4788 => x"a7",
          4789 => x"34",
          4790 => x"33",
          4791 => x"06",
          4792 => x"22",
          4793 => x"33",
          4794 => x"11",
          4795 => x"55",
          4796 => x"90",
          4797 => x"b6",
          4798 => x"18",
          4799 => x"06",
          4800 => x"78",
          4801 => x"38",
          4802 => x"33",
          4803 => x"ea",
          4804 => x"53",
          4805 => x"95",
          4806 => x"db",
          4807 => x"80",
          4808 => x"84",
          4809 => x"57",
          4810 => x"80",
          4811 => x"0b",
          4812 => x"0c",
          4813 => x"04",
          4814 => x"97",
          4815 => x"24",
          4816 => x"75",
          4817 => x"81",
          4818 => x"38",
          4819 => x"51",
          4820 => x"80",
          4821 => x"95",
          4822 => x"39",
          4823 => x"15",
          4824 => x"b6",
          4825 => x"74",
          4826 => x"2e",
          4827 => x"fe",
          4828 => x"53",
          4829 => x"51",
          4830 => x"81",
          4831 => x"ff",
          4832 => x"72",
          4833 => x"91",
          4834 => x"a0",
          4835 => x"3f",
          4836 => x"81",
          4837 => x"54",
          4838 => x"d8",
          4839 => x"39",
          4840 => x"95",
          4841 => x"39",
          4842 => x"51",
          4843 => x"80",
          4844 => x"e4",
          4845 => x"0d",
          4846 => x"ff",
          4847 => x"06",
          4848 => x"83",
          4849 => x"70",
          4850 => x"55",
          4851 => x"73",
          4852 => x"53",
          4853 => x"95",
          4854 => x"a0",
          4855 => x"3f",
          4856 => x"33",
          4857 => x"06",
          4858 => x"53",
          4859 => x"38",
          4860 => x"83",
          4861 => x"fe",
          4862 => x"0b",
          4863 => x"34",
          4864 => x"51",
          4865 => x"fe",
          4866 => x"52",
          4867 => x"d8",
          4868 => x"39",
          4869 => x"02",
          4870 => x"33",
          4871 => x"08",
          4872 => x"81",
          4873 => x"38",
          4874 => x"83",
          4875 => x"8a",
          4876 => x"38",
          4877 => x"82",
          4878 => x"88",
          4879 => x"38",
          4880 => x"88",
          4881 => x"b6",
          4882 => x"f8",
          4883 => x"f8",
          4884 => x"72",
          4885 => x"5e",
          4886 => x"e0",
          4887 => x"a7",
          4888 => x"34",
          4889 => x"33",
          4890 => x"33",
          4891 => x"22",
          4892 => x"12",
          4893 => x"40",
          4894 => x"96",
          4895 => x"f8",
          4896 => x"71",
          4897 => x"40",
          4898 => x"90",
          4899 => x"a7",
          4900 => x"34",
          4901 => x"33",
          4902 => x"06",
          4903 => x"22",
          4904 => x"33",
          4905 => x"11",
          4906 => x"58",
          4907 => x"90",
          4908 => x"b6",
          4909 => x"1d",
          4910 => x"06",
          4911 => x"61",
          4912 => x"38",
          4913 => x"33",
          4914 => x"f1",
          4915 => x"56",
          4916 => x"95",
          4917 => x"84",
          4918 => x"9c",
          4919 => x"78",
          4920 => x"8a",
          4921 => x"25",
          4922 => x"78",
          4923 => x"b3",
          4924 => x"db",
          4925 => x"38",
          4926 => x"b7",
          4927 => x"b6",
          4928 => x"f8",
          4929 => x"f8",
          4930 => x"72",
          4931 => x"40",
          4932 => x"e0",
          4933 => x"a7",
          4934 => x"34",
          4935 => x"33",
          4936 => x"33",
          4937 => x"22",
          4938 => x"12",
          4939 => x"56",
          4940 => x"96",
          4941 => x"f8",
          4942 => x"71",
          4943 => x"57",
          4944 => x"33",
          4945 => x"80",
          4946 => x"b6",
          4947 => x"81",
          4948 => x"f8",
          4949 => x"f8",
          4950 => x"72",
          4951 => x"42",
          4952 => x"83",
          4953 => x"60",
          4954 => x"05",
          4955 => x"58",
          4956 => x"06",
          4957 => x"27",
          4958 => x"77",
          4959 => x"34",
          4960 => x"b8",
          4961 => x"3d",
          4962 => x"9b",
          4963 => x"38",
          4964 => x"83",
          4965 => x"8d",
          4966 => x"06",
          4967 => x"80",
          4968 => x"95",
          4969 => x"84",
          4970 => x"9c",
          4971 => x"78",
          4972 => x"aa",
          4973 => x"56",
          4974 => x"84",
          4975 => x"b7",
          4976 => x"11",
          4977 => x"84",
          4978 => x"78",
          4979 => x"18",
          4980 => x"ff",
          4981 => x"0b",
          4982 => x"1a",
          4983 => x"84",
          4984 => x"9c",
          4985 => x"78",
          4986 => x"e9",
          4987 => x"84",
          4988 => x"84",
          4989 => x"83",
          4990 => x"83",
          4991 => x"72",
          4992 => x"5e",
          4993 => x"b6",
          4994 => x"86",
          4995 => x"1d",
          4996 => x"d8",
          4997 => x"95",
          4998 => x"92",
          4999 => x"29",
          5000 => x"59",
          5001 => x"f8",
          5002 => x"83",
          5003 => x"76",
          5004 => x"5b",
          5005 => x"90",
          5006 => x"b0",
          5007 => x"84",
          5008 => x"70",
          5009 => x"83",
          5010 => x"83",
          5011 => x"72",
          5012 => x"44",
          5013 => x"59",
          5014 => x"33",
          5015 => x"b6",
          5016 => x"1f",
          5017 => x"39",
          5018 => x"51",
          5019 => x"80",
          5020 => x"95",
          5021 => x"39",
          5022 => x"33",
          5023 => x"33",
          5024 => x"06",
          5025 => x"33",
          5026 => x"12",
          5027 => x"80",
          5028 => x"92",
          5029 => x"5d",
          5030 => x"05",
          5031 => x"ff",
          5032 => x"ea",
          5033 => x"59",
          5034 => x"81",
          5035 => x"38",
          5036 => x"06",
          5037 => x"57",
          5038 => x"38",
          5039 => x"83",
          5040 => x"fc",
          5041 => x"0b",
          5042 => x"34",
          5043 => x"b7",
          5044 => x"0b",
          5045 => x"34",
          5046 => x"b7",
          5047 => x"0b",
          5048 => x"0c",
          5049 => x"b8",
          5050 => x"3d",
          5051 => x"f8",
          5052 => x"b8",
          5053 => x"f8",
          5054 => x"b8",
          5055 => x"f8",
          5056 => x"b8",
          5057 => x"0b",
          5058 => x"0c",
          5059 => x"b8",
          5060 => x"3d",
          5061 => x"80",
          5062 => x"81",
          5063 => x"38",
          5064 => x"33",
          5065 => x"33",
          5066 => x"06",
          5067 => x"33",
          5068 => x"06",
          5069 => x"11",
          5070 => x"80",
          5071 => x"92",
          5072 => x"72",
          5073 => x"70",
          5074 => x"06",
          5075 => x"33",
          5076 => x"5c",
          5077 => x"7d",
          5078 => x"fe",
          5079 => x"ff",
          5080 => x"58",
          5081 => x"38",
          5082 => x"83",
          5083 => x"7b",
          5084 => x"7a",
          5085 => x"78",
          5086 => x"72",
          5087 => x"5f",
          5088 => x"b7",
          5089 => x"a7",
          5090 => x"34",
          5091 => x"33",
          5092 => x"33",
          5093 => x"22",
          5094 => x"12",
          5095 => x"40",
          5096 => x"f8",
          5097 => x"83",
          5098 => x"60",
          5099 => x"05",
          5100 => x"f8",
          5101 => x"a7",
          5102 => x"34",
          5103 => x"33",
          5104 => x"06",
          5105 => x"22",
          5106 => x"33",
          5107 => x"11",
          5108 => x"5e",
          5109 => x"90",
          5110 => x"97",
          5111 => x"81",
          5112 => x"ff",
          5113 => x"7c",
          5114 => x"ea",
          5115 => x"d9",
          5116 => x"96",
          5117 => x"19",
          5118 => x"f8",
          5119 => x"f8",
          5120 => x"81",
          5121 => x"ff",
          5122 => x"ac",
          5123 => x"2e",
          5124 => x"78",
          5125 => x"d7",
          5126 => x"2e",
          5127 => x"84",
          5128 => x"5f",
          5129 => x"38",
          5130 => x"56",
          5131 => x"84",
          5132 => x"10",
          5133 => x"c0",
          5134 => x"08",
          5135 => x"83",
          5136 => x"80",
          5137 => x"e7",
          5138 => x"0b",
          5139 => x"0c",
          5140 => x"04",
          5141 => x"33",
          5142 => x"33",
          5143 => x"06",
          5144 => x"33",
          5145 => x"06",
          5146 => x"11",
          5147 => x"80",
          5148 => x"92",
          5149 => x"72",
          5150 => x"70",
          5151 => x"06",
          5152 => x"33",
          5153 => x"5c",
          5154 => x"7f",
          5155 => x"ef",
          5156 => x"7a",
          5157 => x"7a",
          5158 => x"7a",
          5159 => x"72",
          5160 => x"5c",
          5161 => x"b7",
          5162 => x"a7",
          5163 => x"34",
          5164 => x"33",
          5165 => x"33",
          5166 => x"22",
          5167 => x"12",
          5168 => x"56",
          5169 => x"f8",
          5170 => x"83",
          5171 => x"76",
          5172 => x"5a",
          5173 => x"90",
          5174 => x"b0",
          5175 => x"84",
          5176 => x"70",
          5177 => x"83",
          5178 => x"83",
          5179 => x"72",
          5180 => x"5b",
          5181 => x"59",
          5182 => x"33",
          5183 => x"18",
          5184 => x"05",
          5185 => x"06",
          5186 => x"7a",
          5187 => x"38",
          5188 => x"33",
          5189 => x"fb",
          5190 => x"56",
          5191 => x"95",
          5192 => x"70",
          5193 => x"5d",
          5194 => x"26",
          5195 => x"83",
          5196 => x"84",
          5197 => x"83",
          5198 => x"72",
          5199 => x"72",
          5200 => x"72",
          5201 => x"72",
          5202 => x"54",
          5203 => x"5b",
          5204 => x"80",
          5205 => x"a0",
          5206 => x"84",
          5207 => x"83",
          5208 => x"83",
          5209 => x"72",
          5210 => x"5e",
          5211 => x"a0",
          5212 => x"96",
          5213 => x"f8",
          5214 => x"71",
          5215 => x"5e",
          5216 => x"33",
          5217 => x"80",
          5218 => x"b6",
          5219 => x"81",
          5220 => x"f8",
          5221 => x"f8",
          5222 => x"72",
          5223 => x"44",
          5224 => x"83",
          5225 => x"84",
          5226 => x"34",
          5227 => x"70",
          5228 => x"5b",
          5229 => x"27",
          5230 => x"77",
          5231 => x"34",
          5232 => x"82",
          5233 => x"e0",
          5234 => x"84",
          5235 => x"9c",
          5236 => x"83",
          5237 => x"33",
          5238 => x"e0",
          5239 => x"34",
          5240 => x"33",
          5241 => x"06",
          5242 => x"56",
          5243 => x"81",
          5244 => x"e6",
          5245 => x"84",
          5246 => x"9c",
          5247 => x"83",
          5248 => x"33",
          5249 => x"e0",
          5250 => x"34",
          5251 => x"33",
          5252 => x"33",
          5253 => x"33",
          5254 => x"80",
          5255 => x"39",
          5256 => x"42",
          5257 => x"11",
          5258 => x"51",
          5259 => x"3f",
          5260 => x"08",
          5261 => x"f0",
          5262 => x"e5",
          5263 => x"57",
          5264 => x"b7",
          5265 => x"10",
          5266 => x"41",
          5267 => x"05",
          5268 => x"b8",
          5269 => x"fb",
          5270 => x"f8",
          5271 => x"5c",
          5272 => x"1c",
          5273 => x"83",
          5274 => x"84",
          5275 => x"83",
          5276 => x"5b",
          5277 => x"e5",
          5278 => x"d8",
          5279 => x"94",
          5280 => x"95",
          5281 => x"29",
          5282 => x"5b",
          5283 => x"19",
          5284 => x"a7",
          5285 => x"34",
          5286 => x"33",
          5287 => x"33",
          5288 => x"22",
          5289 => x"12",
          5290 => x"56",
          5291 => x"96",
          5292 => x"f8",
          5293 => x"71",
          5294 => x"5e",
          5295 => x"33",
          5296 => x"b0",
          5297 => x"84",
          5298 => x"70",
          5299 => x"83",
          5300 => x"83",
          5301 => x"72",
          5302 => x"41",
          5303 => x"5a",
          5304 => x"33",
          5305 => x"1e",
          5306 => x"70",
          5307 => x"5c",
          5308 => x"26",
          5309 => x"84",
          5310 => x"58",
          5311 => x"38",
          5312 => x"75",
          5313 => x"34",
          5314 => x"b7",
          5315 => x"b6",
          5316 => x"7f",
          5317 => x"bd",
          5318 => x"dc",
          5319 => x"f3",
          5320 => x"52",
          5321 => x"e4",
          5322 => x"84",
          5323 => x"9c",
          5324 => x"84",
          5325 => x"83",
          5326 => x"84",
          5327 => x"83",
          5328 => x"84",
          5329 => x"57",
          5330 => x"92",
          5331 => x"39",
          5332 => x"33",
          5333 => x"34",
          5334 => x"33",
          5335 => x"34",
          5336 => x"33",
          5337 => x"34",
          5338 => x"84",
          5339 => x"5b",
          5340 => x"ff",
          5341 => x"b8",
          5342 => x"7c",
          5343 => x"81",
          5344 => x"38",
          5345 => x"33",
          5346 => x"83",
          5347 => x"81",
          5348 => x"53",
          5349 => x"52",
          5350 => x"52",
          5351 => x"89",
          5352 => x"fe",
          5353 => x"84",
          5354 => x"81",
          5355 => x"f6",
          5356 => x"76",
          5357 => x"a0",
          5358 => x"38",
          5359 => x"f6",
          5360 => x"fd",
          5361 => x"c0",
          5362 => x"84",
          5363 => x"5b",
          5364 => x"ff",
          5365 => x"7b",
          5366 => x"38",
          5367 => x"b8",
          5368 => x"11",
          5369 => x"75",
          5370 => x"a5",
          5371 => x"10",
          5372 => x"05",
          5373 => x"04",
          5374 => x"33",
          5375 => x"2e",
          5376 => x"83",
          5377 => x"84",
          5378 => x"71",
          5379 => x"09",
          5380 => x"72",
          5381 => x"59",
          5382 => x"83",
          5383 => x"fd",
          5384 => x"b7",
          5385 => x"75",
          5386 => x"e7",
          5387 => x"b9",
          5388 => x"70",
          5389 => x"84",
          5390 => x"5d",
          5391 => x"7b",
          5392 => x"38",
          5393 => x"95",
          5394 => x"39",
          5395 => x"f8",
          5396 => x"f8",
          5397 => x"81",
          5398 => x"57",
          5399 => x"fd",
          5400 => x"17",
          5401 => x"f8",
          5402 => x"9c",
          5403 => x"83",
          5404 => x"83",
          5405 => x"84",
          5406 => x"ff",
          5407 => x"76",
          5408 => x"84",
          5409 => x"56",
          5410 => x"94",
          5411 => x"39",
          5412 => x"33",
          5413 => x"2e",
          5414 => x"83",
          5415 => x"84",
          5416 => x"71",
          5417 => x"09",
          5418 => x"72",
          5419 => x"59",
          5420 => x"83",
          5421 => x"fc",
          5422 => x"b7",
          5423 => x"7a",
          5424 => x"c4",
          5425 => x"b8",
          5426 => x"99",
          5427 => x"06",
          5428 => x"84",
          5429 => x"83",
          5430 => x"83",
          5431 => x"72",
          5432 => x"86",
          5433 => x"11",
          5434 => x"22",
          5435 => x"58",
          5436 => x"05",
          5437 => x"ff",
          5438 => x"e8",
          5439 => x"fe",
          5440 => x"5a",
          5441 => x"84",
          5442 => x"92",
          5443 => x"0b",
          5444 => x"34",
          5445 => x"84",
          5446 => x"5a",
          5447 => x"fb",
          5448 => x"b8",
          5449 => x"77",
          5450 => x"81",
          5451 => x"38",
          5452 => x"f6",
          5453 => x"d0",
          5454 => x"e5",
          5455 => x"80",
          5456 => x"38",
          5457 => x"33",
          5458 => x"33",
          5459 => x"84",
          5460 => x"ff",
          5461 => x"56",
          5462 => x"83",
          5463 => x"76",
          5464 => x"34",
          5465 => x"84",
          5466 => x"57",
          5467 => x"8c",
          5468 => x"b8",
          5469 => x"f8",
          5470 => x"61",
          5471 => x"d7",
          5472 => x"59",
          5473 => x"60",
          5474 => x"75",
          5475 => x"f8",
          5476 => x"f4",
          5477 => x"ac",
          5478 => x"ed",
          5479 => x"84",
          5480 => x"57",
          5481 => x"27",
          5482 => x"76",
          5483 => x"b8",
          5484 => x"53",
          5485 => x"8c",
          5486 => x"cd",
          5487 => x"70",
          5488 => x"84",
          5489 => x"58",
          5490 => x"39",
          5491 => x"b7",
          5492 => x"57",
          5493 => x"8d",
          5494 => x"b8",
          5495 => x"83",
          5496 => x"75",
          5497 => x"76",
          5498 => x"51",
          5499 => x"fa",
          5500 => x"b7",
          5501 => x"81",
          5502 => x"b7",
          5503 => x"bb",
          5504 => x"70",
          5505 => x"84",
          5506 => x"ff",
          5507 => x"ff",
          5508 => x"d7",
          5509 => x"ff",
          5510 => x"40",
          5511 => x"59",
          5512 => x"7e",
          5513 => x"77",
          5514 => x"f8",
          5515 => x"81",
          5516 => x"18",
          5517 => x"7f",
          5518 => x"77",
          5519 => x"f8",
          5520 => x"b6",
          5521 => x"11",
          5522 => x"60",
          5523 => x"38",
          5524 => x"83",
          5525 => x"f9",
          5526 => x"b7",
          5527 => x"7e",
          5528 => x"ef",
          5529 => x"b9",
          5530 => x"d7",
          5531 => x"7a",
          5532 => x"94",
          5533 => x"94",
          5534 => x"d8",
          5535 => x"ff",
          5536 => x"95",
          5537 => x"29",
          5538 => x"a0",
          5539 => x"f8",
          5540 => x"40",
          5541 => x"05",
          5542 => x"ff",
          5543 => x"ea",
          5544 => x"59",
          5545 => x"60",
          5546 => x"f0",
          5547 => x"ff",
          5548 => x"7c",
          5549 => x"80",
          5550 => x"fe",
          5551 => x"d7",
          5552 => x"76",
          5553 => x"38",
          5554 => x"75",
          5555 => x"23",
          5556 => x"06",
          5557 => x"41",
          5558 => x"24",
          5559 => x"84",
          5560 => x"56",
          5561 => x"8d",
          5562 => x"16",
          5563 => x"f8",
          5564 => x"81",
          5565 => x"f8",
          5566 => x"57",
          5567 => x"76",
          5568 => x"75",
          5569 => x"05",
          5570 => x"06",
          5571 => x"5c",
          5572 => x"58",
          5573 => x"80",
          5574 => x"b0",
          5575 => x"ff",
          5576 => x"ff",
          5577 => x"29",
          5578 => x"42",
          5579 => x"27",
          5580 => x"84",
          5581 => x"57",
          5582 => x"33",
          5583 => x"e0",
          5584 => x"70",
          5585 => x"34",
          5586 => x"05",
          5587 => x"70",
          5588 => x"34",
          5589 => x"b6",
          5590 => x"b6",
          5591 => x"71",
          5592 => x"40",
          5593 => x"60",
          5594 => x"38",
          5595 => x"33",
          5596 => x"e0",
          5597 => x"70",
          5598 => x"34",
          5599 => x"05",
          5600 => x"70",
          5601 => x"34",
          5602 => x"b6",
          5603 => x"b6",
          5604 => x"71",
          5605 => x"40",
          5606 => x"78",
          5607 => x"38",
          5608 => x"84",
          5609 => x"56",
          5610 => x"87",
          5611 => x"52",
          5612 => x"33",
          5613 => x"3f",
          5614 => x"80",
          5615 => x"d8",
          5616 => x"84",
          5617 => x"5d",
          5618 => x"79",
          5619 => x"38",
          5620 => x"22",
          5621 => x"2e",
          5622 => x"8b",
          5623 => x"f8",
          5624 => x"76",
          5625 => x"83",
          5626 => x"79",
          5627 => x"76",
          5628 => x"ed",
          5629 => x"d7",
          5630 => x"60",
          5631 => x"38",
          5632 => x"06",
          5633 => x"26",
          5634 => x"7b",
          5635 => x"7d",
          5636 => x"76",
          5637 => x"7a",
          5638 => x"70",
          5639 => x"05",
          5640 => x"80",
          5641 => x"5d",
          5642 => x"b0",
          5643 => x"83",
          5644 => x"5d",
          5645 => x"38",
          5646 => x"57",
          5647 => x"38",
          5648 => x"33",
          5649 => x"71",
          5650 => x"71",
          5651 => x"71",
          5652 => x"59",
          5653 => x"77",
          5654 => x"38",
          5655 => x"84",
          5656 => x"7d",
          5657 => x"05",
          5658 => x"77",
          5659 => x"84",
          5660 => x"84",
          5661 => x"41",
          5662 => x"ff",
          5663 => x"ff",
          5664 => x"92",
          5665 => x"29",
          5666 => x"59",
          5667 => x"77",
          5668 => x"76",
          5669 => x"70",
          5670 => x"05",
          5671 => x"76",
          5672 => x"76",
          5673 => x"e0",
          5674 => x"90",
          5675 => x"b6",
          5676 => x"a0",
          5677 => x"19",
          5678 => x"70",
          5679 => x"34",
          5680 => x"76",
          5681 => x"c0",
          5682 => x"e0",
          5683 => x"79",
          5684 => x"05",
          5685 => x"17",
          5686 => x"27",
          5687 => x"a8",
          5688 => x"70",
          5689 => x"5d",
          5690 => x"39",
          5691 => x"33",
          5692 => x"06",
          5693 => x"80",
          5694 => x"84",
          5695 => x"5d",
          5696 => x"f0",
          5697 => x"06",
          5698 => x"f2",
          5699 => x"90",
          5700 => x"70",
          5701 => x"59",
          5702 => x"39",
          5703 => x"17",
          5704 => x"b6",
          5705 => x"7c",
          5706 => x"94",
          5707 => x"d8",
          5708 => x"92",
          5709 => x"d7",
          5710 => x"5f",
          5711 => x"39",
          5712 => x"33",
          5713 => x"75",
          5714 => x"34",
          5715 => x"81",
          5716 => x"56",
          5717 => x"83",
          5718 => x"81",
          5719 => x"07",
          5720 => x"f8",
          5721 => x"39",
          5722 => x"33",
          5723 => x"83",
          5724 => x"83",
          5725 => x"d4",
          5726 => x"90",
          5727 => x"06",
          5728 => x"75",
          5729 => x"34",
          5730 => x"f8",
          5731 => x"9f",
          5732 => x"56",
          5733 => x"90",
          5734 => x"39",
          5735 => x"83",
          5736 => x"81",
          5737 => x"ff",
          5738 => x"f4",
          5739 => x"f8",
          5740 => x"8f",
          5741 => x"83",
          5742 => x"ff",
          5743 => x"f8",
          5744 => x"9f",
          5745 => x"56",
          5746 => x"90",
          5747 => x"39",
          5748 => x"33",
          5749 => x"80",
          5750 => x"75",
          5751 => x"34",
          5752 => x"83",
          5753 => x"81",
          5754 => x"c0",
          5755 => x"83",
          5756 => x"fe",
          5757 => x"f8",
          5758 => x"af",
          5759 => x"56",
          5760 => x"90",
          5761 => x"39",
          5762 => x"33",
          5763 => x"86",
          5764 => x"83",
          5765 => x"fe",
          5766 => x"f8",
          5767 => x"fc",
          5768 => x"56",
          5769 => x"90",
          5770 => x"39",
          5771 => x"33",
          5772 => x"82",
          5773 => x"83",
          5774 => x"fe",
          5775 => x"f8",
          5776 => x"f8",
          5777 => x"83",
          5778 => x"fd",
          5779 => x"f8",
          5780 => x"f0",
          5781 => x"83",
          5782 => x"fd",
          5783 => x"f8",
          5784 => x"f0",
          5785 => x"83",
          5786 => x"fd",
          5787 => x"f8",
          5788 => x"df",
          5789 => x"07",
          5790 => x"f8",
          5791 => x"cc",
          5792 => x"90",
          5793 => x"06",
          5794 => x"75",
          5795 => x"34",
          5796 => x"80",
          5797 => x"95",
          5798 => x"81",
          5799 => x"3f",
          5800 => x"84",
          5801 => x"83",
          5802 => x"84",
          5803 => x"83",
          5804 => x"84",
          5805 => x"59",
          5806 => x"92",
          5807 => x"84",
          5808 => x"e8",
          5809 => x"0b",
          5810 => x"34",
          5811 => x"b8",
          5812 => x"3d",
          5813 => x"83",
          5814 => x"83",
          5815 => x"70",
          5816 => x"58",
          5817 => x"e7",
          5818 => x"b7",
          5819 => x"3d",
          5820 => x"d8",
          5821 => x"f9",
          5822 => x"b8",
          5823 => x"38",
          5824 => x"08",
          5825 => x"0c",
          5826 => x"b7",
          5827 => x"0b",
          5828 => x"0c",
          5829 => x"04",
          5830 => x"95",
          5831 => x"39",
          5832 => x"33",
          5833 => x"5c",
          5834 => x"e5",
          5835 => x"83",
          5836 => x"02",
          5837 => x"22",
          5838 => x"1e",
          5839 => x"84",
          5840 => x"ca",
          5841 => x"83",
          5842 => x"80",
          5843 => x"d1",
          5844 => x"f8",
          5845 => x"81",
          5846 => x"ff",
          5847 => x"d8",
          5848 => x"83",
          5849 => x"80",
          5850 => x"d0",
          5851 => x"98",
          5852 => x"fe",
          5853 => x"ef",
          5854 => x"f8",
          5855 => x"05",
          5856 => x"9f",
          5857 => x"58",
          5858 => x"a6",
          5859 => x"81",
          5860 => x"84",
          5861 => x"40",
          5862 => x"ee",
          5863 => x"83",
          5864 => x"ee",
          5865 => x"f8",
          5866 => x"05",
          5867 => x"9f",
          5868 => x"58",
          5869 => x"e2",
          5870 => x"94",
          5871 => x"84",
          5872 => x"ff",
          5873 => x"56",
          5874 => x"f3",
          5875 => x"57",
          5876 => x"84",
          5877 => x"70",
          5878 => x"58",
          5879 => x"26",
          5880 => x"83",
          5881 => x"84",
          5882 => x"70",
          5883 => x"83",
          5884 => x"71",
          5885 => x"86",
          5886 => x"05",
          5887 => x"22",
          5888 => x"7e",
          5889 => x"83",
          5890 => x"83",
          5891 => x"5d",
          5892 => x"5f",
          5893 => x"2e",
          5894 => x"79",
          5895 => x"06",
          5896 => x"57",
          5897 => x"84",
          5898 => x"b6",
          5899 => x"76",
          5900 => x"98",
          5901 => x"56",
          5902 => x"92",
          5903 => x"ff",
          5904 => x"57",
          5905 => x"24",
          5906 => x"84",
          5907 => x"56",
          5908 => x"82",
          5909 => x"16",
          5910 => x"f8",
          5911 => x"81",
          5912 => x"f8",
          5913 => x"57",
          5914 => x"76",
          5915 => x"75",
          5916 => x"05",
          5917 => x"06",
          5918 => x"5c",
          5919 => x"58",
          5920 => x"80",
          5921 => x"b0",
          5922 => x"ff",
          5923 => x"ff",
          5924 => x"29",
          5925 => x"42",
          5926 => x"27",
          5927 => x"84",
          5928 => x"57",
          5929 => x"33",
          5930 => x"e0",
          5931 => x"70",
          5932 => x"34",
          5933 => x"05",
          5934 => x"70",
          5935 => x"34",
          5936 => x"b6",
          5937 => x"b6",
          5938 => x"71",
          5939 => x"41",
          5940 => x"76",
          5941 => x"38",
          5942 => x"33",
          5943 => x"e0",
          5944 => x"70",
          5945 => x"34",
          5946 => x"05",
          5947 => x"70",
          5948 => x"34",
          5949 => x"b6",
          5950 => x"b6",
          5951 => x"71",
          5952 => x"41",
          5953 => x"78",
          5954 => x"38",
          5955 => x"83",
          5956 => x"33",
          5957 => x"e0",
          5958 => x"34",
          5959 => x"33",
          5960 => x"33",
          5961 => x"22",
          5962 => x"33",
          5963 => x"5d",
          5964 => x"76",
          5965 => x"84",
          5966 => x"70",
          5967 => x"ff",
          5968 => x"58",
          5969 => x"83",
          5970 => x"79",
          5971 => x"23",
          5972 => x"06",
          5973 => x"5a",
          5974 => x"83",
          5975 => x"76",
          5976 => x"34",
          5977 => x"33",
          5978 => x"06",
          5979 => x"59",
          5980 => x"27",
          5981 => x"80",
          5982 => x"f8",
          5983 => x"88",
          5984 => x"95",
          5985 => x"84",
          5986 => x"ff",
          5987 => x"56",
          5988 => x"ef",
          5989 => x"57",
          5990 => x"75",
          5991 => x"81",
          5992 => x"38",
          5993 => x"33",
          5994 => x"06",
          5995 => x"33",
          5996 => x"5d",
          5997 => x"2e",
          5998 => x"f4",
          5999 => x"a1",
          6000 => x"56",
          6001 => x"94",
          6002 => x"39",
          6003 => x"75",
          6004 => x"23",
          6005 => x"7c",
          6006 => x"75",
          6007 => x"34",
          6008 => x"77",
          6009 => x"77",
          6010 => x"8d",
          6011 => x"70",
          6012 => x"34",
          6013 => x"33",
          6014 => x"05",
          6015 => x"7a",
          6016 => x"38",
          6017 => x"81",
          6018 => x"83",
          6019 => x"77",
          6020 => x"59",
          6021 => x"27",
          6022 => x"d3",
          6023 => x"31",
          6024 => x"f8",
          6025 => x"a8",
          6026 => x"83",
          6027 => x"fc",
          6028 => x"83",
          6029 => x"fc",
          6030 => x"0b",
          6031 => x"23",
          6032 => x"80",
          6033 => x"94",
          6034 => x"39",
          6035 => x"18",
          6036 => x"b6",
          6037 => x"77",
          6038 => x"83",
          6039 => x"e9",
          6040 => x"3d",
          6041 => x"05",
          6042 => x"da",
          6043 => x"72",
          6044 => x"38",
          6045 => x"9c",
          6046 => x"84",
          6047 => x"85",
          6048 => x"76",
          6049 => x"d7",
          6050 => x"0b",
          6051 => x"0c",
          6052 => x"04",
          6053 => x"02",
          6054 => x"5c",
          6055 => x"f6",
          6056 => x"81",
          6057 => x"f6",
          6058 => x"58",
          6059 => x"74",
          6060 => x"d6",
          6061 => x"56",
          6062 => x"e8",
          6063 => x"78",
          6064 => x"0c",
          6065 => x"04",
          6066 => x"08",
          6067 => x"73",
          6068 => x"38",
          6069 => x"70",
          6070 => x"70",
          6071 => x"2a",
          6072 => x"58",
          6073 => x"c4",
          6074 => x"80",
          6075 => x"2e",
          6076 => x"83",
          6077 => x"7b",
          6078 => x"30",
          6079 => x"76",
          6080 => x"5d",
          6081 => x"85",
          6082 => x"b6",
          6083 => x"f8",
          6084 => x"f8",
          6085 => x"71",
          6086 => x"a7",
          6087 => x"83",
          6088 => x"5b",
          6089 => x"79",
          6090 => x"83",
          6091 => x"83",
          6092 => x"58",
          6093 => x"74",
          6094 => x"8c",
          6095 => x"54",
          6096 => x"80",
          6097 => x"0b",
          6098 => x"88",
          6099 => x"98",
          6100 => x"75",
          6101 => x"38",
          6102 => x"84",
          6103 => x"83",
          6104 => x"34",
          6105 => x"81",
          6106 => x"55",
          6107 => x"27",
          6108 => x"54",
          6109 => x"14",
          6110 => x"ff",
          6111 => x"8e",
          6112 => x"54",
          6113 => x"2e",
          6114 => x"72",
          6115 => x"86",
          6116 => x"83",
          6117 => x"34",
          6118 => x"06",
          6119 => x"ff",
          6120 => x"38",
          6121 => x"a2",
          6122 => x"f6",
          6123 => x"83",
          6124 => x"34",
          6125 => x"81",
          6126 => x"5e",
          6127 => x"ff",
          6128 => x"f6",
          6129 => x"98",
          6130 => x"25",
          6131 => x"75",
          6132 => x"34",
          6133 => x"06",
          6134 => x"81",
          6135 => x"06",
          6136 => x"72",
          6137 => x"e7",
          6138 => x"83",
          6139 => x"73",
          6140 => x"53",
          6141 => x"85",
          6142 => x"0b",
          6143 => x"34",
          6144 => x"f6",
          6145 => x"f6",
          6146 => x"f6",
          6147 => x"83",
          6148 => x"83",
          6149 => x"5d",
          6150 => x"5c",
          6151 => x"f6",
          6152 => x"55",
          6153 => x"2e",
          6154 => x"f6",
          6155 => x"54",
          6156 => x"82",
          6157 => x"f6",
          6158 => x"53",
          6159 => x"2e",
          6160 => x"f6",
          6161 => x"54",
          6162 => x"38",
          6163 => x"06",
          6164 => x"ff",
          6165 => x"83",
          6166 => x"33",
          6167 => x"2e",
          6168 => x"74",
          6169 => x"53",
          6170 => x"2e",
          6171 => x"83",
          6172 => x"33",
          6173 => x"27",
          6174 => x"83",
          6175 => x"87",
          6176 => x"c0",
          6177 => x"54",
          6178 => x"27",
          6179 => x"81",
          6180 => x"98",
          6181 => x"f6",
          6182 => x"81",
          6183 => x"ff",
          6184 => x"89",
          6185 => x"f6",
          6186 => x"f6",
          6187 => x"83",
          6188 => x"fe",
          6189 => x"72",
          6190 => x"8b",
          6191 => x"10",
          6192 => x"05",
          6193 => x"04",
          6194 => x"08",
          6195 => x"2e",
          6196 => x"f4",
          6197 => x"98",
          6198 => x"5e",
          6199 => x"fc",
          6200 => x"0b",
          6201 => x"33",
          6202 => x"81",
          6203 => x"74",
          6204 => x"f6",
          6205 => x"c0",
          6206 => x"83",
          6207 => x"73",
          6208 => x"58",
          6209 => x"94",
          6210 => x"96",
          6211 => x"84",
          6212 => x"33",
          6213 => x"f0",
          6214 => x"39",
          6215 => x"08",
          6216 => x"2e",
          6217 => x"72",
          6218 => x"f4",
          6219 => x"76",
          6220 => x"54",
          6221 => x"80",
          6222 => x"39",
          6223 => x"57",
          6224 => x"81",
          6225 => x"79",
          6226 => x"81",
          6227 => x"38",
          6228 => x"80",
          6229 => x"81",
          6230 => x"38",
          6231 => x"06",
          6232 => x"27",
          6233 => x"54",
          6234 => x"25",
          6235 => x"80",
          6236 => x"81",
          6237 => x"ff",
          6238 => x"81",
          6239 => x"72",
          6240 => x"2b",
          6241 => x"58",
          6242 => x"24",
          6243 => x"10",
          6244 => x"10",
          6245 => x"83",
          6246 => x"83",
          6247 => x"70",
          6248 => x"54",
          6249 => x"98",
          6250 => x"f6",
          6251 => x"fd",
          6252 => x"59",
          6253 => x"ff",
          6254 => x"81",
          6255 => x"ff",
          6256 => x"59",
          6257 => x"78",
          6258 => x"9f",
          6259 => x"84",
          6260 => x"54",
          6261 => x"2e",
          6262 => x"7b",
          6263 => x"30",
          6264 => x"76",
          6265 => x"56",
          6266 => x"7b",
          6267 => x"81",
          6268 => x"38",
          6269 => x"f9",
          6270 => x"53",
          6271 => x"10",
          6272 => x"05",
          6273 => x"54",
          6274 => x"83",
          6275 => x"13",
          6276 => x"06",
          6277 => x"73",
          6278 => x"84",
          6279 => x"53",
          6280 => x"f9",
          6281 => x"b6",
          6282 => x"74",
          6283 => x"78",
          6284 => x"52",
          6285 => x"d4",
          6286 => x"b8",
          6287 => x"3d",
          6288 => x"76",
          6289 => x"54",
          6290 => x"72",
          6291 => x"92",
          6292 => x"ac",
          6293 => x"05",
          6294 => x"f6",
          6295 => x"fa",
          6296 => x"0b",
          6297 => x"15",
          6298 => x"83",
          6299 => x"34",
          6300 => x"f6",
          6301 => x"fa",
          6302 => x"81",
          6303 => x"72",
          6304 => x"fc",
          6305 => x"f6",
          6306 => x"55",
          6307 => x"fc",
          6308 => x"81",
          6309 => x"73",
          6310 => x"81",
          6311 => x"38",
          6312 => x"08",
          6313 => x"87",
          6314 => x"08",
          6315 => x"73",
          6316 => x"38",
          6317 => x"9c",
          6318 => x"b8",
          6319 => x"ff",
          6320 => x"d7",
          6321 => x"83",
          6322 => x"34",
          6323 => x"72",
          6324 => x"34",
          6325 => x"06",
          6326 => x"9e",
          6327 => x"f6",
          6328 => x"0b",
          6329 => x"33",
          6330 => x"08",
          6331 => x"33",
          6332 => x"c0",
          6333 => x"bf",
          6334 => x"42",
          6335 => x"56",
          6336 => x"79",
          6337 => x"81",
          6338 => x"38",
          6339 => x"81",
          6340 => x"38",
          6341 => x"09",
          6342 => x"c0",
          6343 => x"39",
          6344 => x"81",
          6345 => x"98",
          6346 => x"84",
          6347 => x"57",
          6348 => x"38",
          6349 => x"84",
          6350 => x"ff",
          6351 => x"39",
          6352 => x"b6",
          6353 => x"54",
          6354 => x"81",
          6355 => x"b6",
          6356 => x"59",
          6357 => x"81",
          6358 => x"c4",
          6359 => x"f7",
          6360 => x"0b",
          6361 => x"0c",
          6362 => x"84",
          6363 => x"70",
          6364 => x"ff",
          6365 => x"54",
          6366 => x"83",
          6367 => x"74",
          6368 => x"23",
          6369 => x"06",
          6370 => x"53",
          6371 => x"83",
          6372 => x"73",
          6373 => x"34",
          6374 => x"33",
          6375 => x"06",
          6376 => x"53",
          6377 => x"83",
          6378 => x"72",
          6379 => x"34",
          6380 => x"b7",
          6381 => x"83",
          6382 => x"a5",
          6383 => x"f6",
          6384 => x"54",
          6385 => x"84",
          6386 => x"83",
          6387 => x"fe",
          6388 => x"81",
          6389 => x"e8",
          6390 => x"c8",
          6391 => x"bb",
          6392 => x"0d",
          6393 => x"ac",
          6394 => x"0d",
          6395 => x"0d",
          6396 => x"f2",
          6397 => x"57",
          6398 => x"33",
          6399 => x"83",
          6400 => x"51",
          6401 => x"34",
          6402 => x"f2",
          6403 => x"56",
          6404 => x"15",
          6405 => x"86",
          6406 => x"34",
          6407 => x"9c",
          6408 => x"f0",
          6409 => x"ce",
          6410 => x"87",
          6411 => x"08",
          6412 => x"98",
          6413 => x"70",
          6414 => x"38",
          6415 => x"87",
          6416 => x"08",
          6417 => x"73",
          6418 => x"71",
          6419 => x"db",
          6420 => x"98",
          6421 => x"ff",
          6422 => x"27",
          6423 => x"71",
          6424 => x"2e",
          6425 => x"87",
          6426 => x"08",
          6427 => x"05",
          6428 => x"98",
          6429 => x"87",
          6430 => x"08",
          6431 => x"2e",
          6432 => x"14",
          6433 => x"98",
          6434 => x"52",
          6435 => x"87",
          6436 => x"ff",
          6437 => x"87",
          6438 => x"08",
          6439 => x"26",
          6440 => x"52",
          6441 => x"16",
          6442 => x"06",
          6443 => x"80",
          6444 => x"74",
          6445 => x"52",
          6446 => x"38",
          6447 => x"8a",
          6448 => x"b8",
          6449 => x"3d",
          6450 => x"0b",
          6451 => x"0c",
          6452 => x"04",
          6453 => x"79",
          6454 => x"a3",
          6455 => x"52",
          6456 => x"f2",
          6457 => x"88",
          6458 => x"80",
          6459 => x"75",
          6460 => x"51",
          6461 => x"71",
          6462 => x"72",
          6463 => x"70",
          6464 => x"71",
          6465 => x"75",
          6466 => x"72",
          6467 => x"83",
          6468 => x"52",
          6469 => x"34",
          6470 => x"08",
          6471 => x"71",
          6472 => x"83",
          6473 => x"55",
          6474 => x"81",
          6475 => x"0b",
          6476 => x"e8",
          6477 => x"98",
          6478 => x"f2",
          6479 => x"80",
          6480 => x"53",
          6481 => x"9c",
          6482 => x"c0",
          6483 => x"51",
          6484 => x"f6",
          6485 => x"33",
          6486 => x"9c",
          6487 => x"74",
          6488 => x"38",
          6489 => x"2e",
          6490 => x"c0",
          6491 => x"51",
          6492 => x"73",
          6493 => x"38",
          6494 => x"ff",
          6495 => x"38",
          6496 => x"9c",
          6497 => x"90",
          6498 => x"c0",
          6499 => x"52",
          6500 => x"9c",
          6501 => x"72",
          6502 => x"81",
          6503 => x"c0",
          6504 => x"52",
          6505 => x"27",
          6506 => x"81",
          6507 => x"38",
          6508 => x"a4",
          6509 => x"75",
          6510 => x"ff",
          6511 => x"ff",
          6512 => x"ff",
          6513 => x"75",
          6514 => x"c7",
          6515 => x"ff",
          6516 => x"fe",
          6517 => x"51",
          6518 => x"06",
          6519 => x"38",
          6520 => x"7b",
          6521 => x"55",
          6522 => x"73",
          6523 => x"71",
          6524 => x"53",
          6525 => x"81",
          6526 => x"72",
          6527 => x"38",
          6528 => x"e4",
          6529 => x"0d",
          6530 => x"84",
          6531 => x"88",
          6532 => x"ff",
          6533 => x"fa",
          6534 => x"02",
          6535 => x"05",
          6536 => x"80",
          6537 => x"f0",
          6538 => x"2b",
          6539 => x"80",
          6540 => x"98",
          6541 => x"55",
          6542 => x"83",
          6543 => x"90",
          6544 => x"84",
          6545 => x"90",
          6546 => x"85",
          6547 => x"86",
          6548 => x"83",
          6549 => x"80",
          6550 => x"80",
          6551 => x"55",
          6552 => x"27",
          6553 => x"70",
          6554 => x"33",
          6555 => x"05",
          6556 => x"71",
          6557 => x"83",
          6558 => x"54",
          6559 => x"34",
          6560 => x"08",
          6561 => x"75",
          6562 => x"83",
          6563 => x"55",
          6564 => x"81",
          6565 => x"0b",
          6566 => x"e8",
          6567 => x"98",
          6568 => x"f2",
          6569 => x"80",
          6570 => x"53",
          6571 => x"9c",
          6572 => x"c0",
          6573 => x"51",
          6574 => x"f6",
          6575 => x"33",
          6576 => x"9c",
          6577 => x"74",
          6578 => x"38",
          6579 => x"2e",
          6580 => x"c0",
          6581 => x"51",
          6582 => x"73",
          6583 => x"38",
          6584 => x"ff",
          6585 => x"38",
          6586 => x"9c",
          6587 => x"90",
          6588 => x"c0",
          6589 => x"52",
          6590 => x"9c",
          6591 => x"72",
          6592 => x"81",
          6593 => x"c0",
          6594 => x"52",
          6595 => x"27",
          6596 => x"81",
          6597 => x"38",
          6598 => x"a4",
          6599 => x"75",
          6600 => x"ff",
          6601 => x"ff",
          6602 => x"ff",
          6603 => x"75",
          6604 => x"38",
          6605 => x"06",
          6606 => x"d5",
          6607 => x"70",
          6608 => x"54",
          6609 => x"83",
          6610 => x"76",
          6611 => x"0c",
          6612 => x"04",
          6613 => x"39",
          6614 => x"83",
          6615 => x"51",
          6616 => x"34",
          6617 => x"f2",
          6618 => x"56",
          6619 => x"16",
          6620 => x"86",
          6621 => x"34",
          6622 => x"9c",
          6623 => x"f0",
          6624 => x"ce",
          6625 => x"87",
          6626 => x"08",
          6627 => x"98",
          6628 => x"72",
          6629 => x"38",
          6630 => x"87",
          6631 => x"08",
          6632 => x"74",
          6633 => x"71",
          6634 => x"db",
          6635 => x"98",
          6636 => x"ff",
          6637 => x"27",
          6638 => x"71",
          6639 => x"2e",
          6640 => x"87",
          6641 => x"08",
          6642 => x"05",
          6643 => x"98",
          6644 => x"87",
          6645 => x"08",
          6646 => x"2e",
          6647 => x"15",
          6648 => x"98",
          6649 => x"52",
          6650 => x"87",
          6651 => x"ff",
          6652 => x"87",
          6653 => x"08",
          6654 => x"26",
          6655 => x"52",
          6656 => x"16",
          6657 => x"06",
          6658 => x"80",
          6659 => x"72",
          6660 => x"54",
          6661 => x"38",
          6662 => x"3d",
          6663 => x"e8",
          6664 => x"d0",
          6665 => x"0d",
          6666 => x"0d",
          6667 => x"08",
          6668 => x"83",
          6669 => x"ff",
          6670 => x"83",
          6671 => x"70",
          6672 => x"33",
          6673 => x"71",
          6674 => x"77",
          6675 => x"81",
          6676 => x"98",
          6677 => x"2b",
          6678 => x"41",
          6679 => x"57",
          6680 => x"57",
          6681 => x"24",
          6682 => x"72",
          6683 => x"33",
          6684 => x"71",
          6685 => x"83",
          6686 => x"05",
          6687 => x"12",
          6688 => x"2b",
          6689 => x"07",
          6690 => x"52",
          6691 => x"80",
          6692 => x"9e",
          6693 => x"33",
          6694 => x"71",
          6695 => x"83",
          6696 => x"05",
          6697 => x"52",
          6698 => x"74",
          6699 => x"73",
          6700 => x"54",
          6701 => x"34",
          6702 => x"08",
          6703 => x"12",
          6704 => x"33",
          6705 => x"07",
          6706 => x"5c",
          6707 => x"51",
          6708 => x"34",
          6709 => x"34",
          6710 => x"08",
          6711 => x"0b",
          6712 => x"80",
          6713 => x"34",
          6714 => x"08",
          6715 => x"14",
          6716 => x"14",
          6717 => x"d4",
          6718 => x"33",
          6719 => x"71",
          6720 => x"82",
          6721 => x"70",
          6722 => x"58",
          6723 => x"72",
          6724 => x"13",
          6725 => x"0d",
          6726 => x"33",
          6727 => x"71",
          6728 => x"83",
          6729 => x"11",
          6730 => x"85",
          6731 => x"88",
          6732 => x"88",
          6733 => x"54",
          6734 => x"58",
          6735 => x"34",
          6736 => x"34",
          6737 => x"08",
          6738 => x"11",
          6739 => x"33",
          6740 => x"71",
          6741 => x"56",
          6742 => x"72",
          6743 => x"33",
          6744 => x"71",
          6745 => x"70",
          6746 => x"55",
          6747 => x"86",
          6748 => x"87",
          6749 => x"b8",
          6750 => x"70",
          6751 => x"33",
          6752 => x"07",
          6753 => x"06",
          6754 => x"5a",
          6755 => x"76",
          6756 => x"81",
          6757 => x"b8",
          6758 => x"17",
          6759 => x"12",
          6760 => x"2b",
          6761 => x"07",
          6762 => x"33",
          6763 => x"71",
          6764 => x"70",
          6765 => x"ff",
          6766 => x"05",
          6767 => x"54",
          6768 => x"5c",
          6769 => x"52",
          6770 => x"34",
          6771 => x"34",
          6772 => x"08",
          6773 => x"33",
          6774 => x"71",
          6775 => x"83",
          6776 => x"05",
          6777 => x"12",
          6778 => x"2b",
          6779 => x"ff",
          6780 => x"2a",
          6781 => x"55",
          6782 => x"52",
          6783 => x"70",
          6784 => x"84",
          6785 => x"70",
          6786 => x"33",
          6787 => x"71",
          6788 => x"83",
          6789 => x"05",
          6790 => x"12",
          6791 => x"2b",
          6792 => x"07",
          6793 => x"52",
          6794 => x"53",
          6795 => x"fc",
          6796 => x"33",
          6797 => x"71",
          6798 => x"82",
          6799 => x"70",
          6800 => x"59",
          6801 => x"34",
          6802 => x"34",
          6803 => x"08",
          6804 => x"33",
          6805 => x"71",
          6806 => x"83",
          6807 => x"05",
          6808 => x"83",
          6809 => x"88",
          6810 => x"88",
          6811 => x"5c",
          6812 => x"52",
          6813 => x"15",
          6814 => x"15",
          6815 => x"0d",
          6816 => x"0d",
          6817 => x"d4",
          6818 => x"76",
          6819 => x"38",
          6820 => x"86",
          6821 => x"fb",
          6822 => x"3d",
          6823 => x"ff",
          6824 => x"b8",
          6825 => x"80",
          6826 => x"d0",
          6827 => x"80",
          6828 => x"84",
          6829 => x"fe",
          6830 => x"84",
          6831 => x"55",
          6832 => x"81",
          6833 => x"34",
          6834 => x"08",
          6835 => x"15",
          6836 => x"85",
          6837 => x"b8",
          6838 => x"76",
          6839 => x"81",
          6840 => x"34",
          6841 => x"08",
          6842 => x"22",
          6843 => x"80",
          6844 => x"83",
          6845 => x"70",
          6846 => x"51",
          6847 => x"88",
          6848 => x"89",
          6849 => x"b8",
          6850 => x"10",
          6851 => x"b8",
          6852 => x"f8",
          6853 => x"76",
          6854 => x"81",
          6855 => x"34",
          6856 => x"f7",
          6857 => x"52",
          6858 => x"51",
          6859 => x"8e",
          6860 => x"83",
          6861 => x"70",
          6862 => x"06",
          6863 => x"83",
          6864 => x"84",
          6865 => x"84",
          6866 => x"12",
          6867 => x"2b",
          6868 => x"59",
          6869 => x"81",
          6870 => x"75",
          6871 => x"cc",
          6872 => x"10",
          6873 => x"33",
          6874 => x"71",
          6875 => x"70",
          6876 => x"06",
          6877 => x"83",
          6878 => x"70",
          6879 => x"53",
          6880 => x"52",
          6881 => x"8a",
          6882 => x"2e",
          6883 => x"73",
          6884 => x"12",
          6885 => x"33",
          6886 => x"07",
          6887 => x"c1",
          6888 => x"ff",
          6889 => x"38",
          6890 => x"56",
          6891 => x"2b",
          6892 => x"33",
          6893 => x"71",
          6894 => x"70",
          6895 => x"06",
          6896 => x"56",
          6897 => x"79",
          6898 => x"81",
          6899 => x"74",
          6900 => x"8d",
          6901 => x"78",
          6902 => x"85",
          6903 => x"2e",
          6904 => x"74",
          6905 => x"2b",
          6906 => x"82",
          6907 => x"70",
          6908 => x"5c",
          6909 => x"76",
          6910 => x"81",
          6911 => x"b8",
          6912 => x"76",
          6913 => x"53",
          6914 => x"34",
          6915 => x"34",
          6916 => x"08",
          6917 => x"33",
          6918 => x"71",
          6919 => x"70",
          6920 => x"ff",
          6921 => x"05",
          6922 => x"ff",
          6923 => x"2a",
          6924 => x"57",
          6925 => x"75",
          6926 => x"72",
          6927 => x"53",
          6928 => x"34",
          6929 => x"08",
          6930 => x"74",
          6931 => x"15",
          6932 => x"d4",
          6933 => x"86",
          6934 => x"12",
          6935 => x"2b",
          6936 => x"07",
          6937 => x"5c",
          6938 => x"75",
          6939 => x"72",
          6940 => x"84",
          6941 => x"70",
          6942 => x"05",
          6943 => x"87",
          6944 => x"88",
          6945 => x"88",
          6946 => x"58",
          6947 => x"15",
          6948 => x"15",
          6949 => x"d4",
          6950 => x"84",
          6951 => x"12",
          6952 => x"2b",
          6953 => x"07",
          6954 => x"5a",
          6955 => x"75",
          6956 => x"72",
          6957 => x"84",
          6958 => x"70",
          6959 => x"05",
          6960 => x"85",
          6961 => x"88",
          6962 => x"88",
          6963 => x"57",
          6964 => x"15",
          6965 => x"15",
          6966 => x"d4",
          6967 => x"05",
          6968 => x"b8",
          6969 => x"3d",
          6970 => x"14",
          6971 => x"33",
          6972 => x"71",
          6973 => x"79",
          6974 => x"33",
          6975 => x"71",
          6976 => x"70",
          6977 => x"5b",
          6978 => x"52",
          6979 => x"34",
          6980 => x"34",
          6981 => x"08",
          6982 => x"11",
          6983 => x"33",
          6984 => x"71",
          6985 => x"74",
          6986 => x"33",
          6987 => x"71",
          6988 => x"70",
          6989 => x"5d",
          6990 => x"5b",
          6991 => x"86",
          6992 => x"87",
          6993 => x"b8",
          6994 => x"70",
          6995 => x"33",
          6996 => x"07",
          6997 => x"06",
          6998 => x"59",
          6999 => x"75",
          7000 => x"81",
          7001 => x"b8",
          7002 => x"84",
          7003 => x"f1",
          7004 => x"0d",
          7005 => x"d4",
          7006 => x"76",
          7007 => x"38",
          7008 => x"8a",
          7009 => x"b8",
          7010 => x"3d",
          7011 => x"51",
          7012 => x"84",
          7013 => x"84",
          7014 => x"89",
          7015 => x"84",
          7016 => x"84",
          7017 => x"a0",
          7018 => x"b8",
          7019 => x"80",
          7020 => x"52",
          7021 => x"51",
          7022 => x"3f",
          7023 => x"08",
          7024 => x"34",
          7025 => x"16",
          7026 => x"d4",
          7027 => x"84",
          7028 => x"0b",
          7029 => x"84",
          7030 => x"56",
          7031 => x"34",
          7032 => x"17",
          7033 => x"d4",
          7034 => x"d0",
          7035 => x"fe",
          7036 => x"70",
          7037 => x"06",
          7038 => x"58",
          7039 => x"74",
          7040 => x"73",
          7041 => x"84",
          7042 => x"70",
          7043 => x"84",
          7044 => x"05",
          7045 => x"55",
          7046 => x"34",
          7047 => x"15",
          7048 => x"77",
          7049 => x"dd",
          7050 => x"39",
          7051 => x"65",
          7052 => x"80",
          7053 => x"d4",
          7054 => x"41",
          7055 => x"84",
          7056 => x"80",
          7057 => x"38",
          7058 => x"88",
          7059 => x"54",
          7060 => x"8f",
          7061 => x"05",
          7062 => x"05",
          7063 => x"ff",
          7064 => x"73",
          7065 => x"06",
          7066 => x"83",
          7067 => x"ff",
          7068 => x"83",
          7069 => x"70",
          7070 => x"33",
          7071 => x"07",
          7072 => x"70",
          7073 => x"06",
          7074 => x"10",
          7075 => x"83",
          7076 => x"70",
          7077 => x"33",
          7078 => x"07",
          7079 => x"70",
          7080 => x"42",
          7081 => x"53",
          7082 => x"5c",
          7083 => x"5e",
          7084 => x"7a",
          7085 => x"38",
          7086 => x"83",
          7087 => x"88",
          7088 => x"10",
          7089 => x"70",
          7090 => x"33",
          7091 => x"71",
          7092 => x"53",
          7093 => x"56",
          7094 => x"24",
          7095 => x"7a",
          7096 => x"f6",
          7097 => x"58",
          7098 => x"87",
          7099 => x"80",
          7100 => x"38",
          7101 => x"77",
          7102 => x"be",
          7103 => x"59",
          7104 => x"92",
          7105 => x"1e",
          7106 => x"12",
          7107 => x"2b",
          7108 => x"07",
          7109 => x"33",
          7110 => x"71",
          7111 => x"90",
          7112 => x"43",
          7113 => x"57",
          7114 => x"60",
          7115 => x"38",
          7116 => x"11",
          7117 => x"33",
          7118 => x"71",
          7119 => x"7a",
          7120 => x"33",
          7121 => x"71",
          7122 => x"83",
          7123 => x"05",
          7124 => x"85",
          7125 => x"88",
          7126 => x"88",
          7127 => x"48",
          7128 => x"58",
          7129 => x"56",
          7130 => x"34",
          7131 => x"34",
          7132 => x"08",
          7133 => x"11",
          7134 => x"33",
          7135 => x"71",
          7136 => x"74",
          7137 => x"33",
          7138 => x"71",
          7139 => x"70",
          7140 => x"42",
          7141 => x"57",
          7142 => x"86",
          7143 => x"87",
          7144 => x"b8",
          7145 => x"70",
          7146 => x"33",
          7147 => x"07",
          7148 => x"06",
          7149 => x"5a",
          7150 => x"76",
          7151 => x"81",
          7152 => x"b8",
          7153 => x"1f",
          7154 => x"83",
          7155 => x"8b",
          7156 => x"2b",
          7157 => x"73",
          7158 => x"33",
          7159 => x"07",
          7160 => x"41",
          7161 => x"5f",
          7162 => x"79",
          7163 => x"81",
          7164 => x"b8",
          7165 => x"1f",
          7166 => x"12",
          7167 => x"2b",
          7168 => x"07",
          7169 => x"14",
          7170 => x"33",
          7171 => x"07",
          7172 => x"41",
          7173 => x"5f",
          7174 => x"79",
          7175 => x"75",
          7176 => x"84",
          7177 => x"70",
          7178 => x"33",
          7179 => x"71",
          7180 => x"66",
          7181 => x"70",
          7182 => x"52",
          7183 => x"05",
          7184 => x"fe",
          7185 => x"84",
          7186 => x"1e",
          7187 => x"65",
          7188 => x"83",
          7189 => x"5d",
          7190 => x"62",
          7191 => x"38",
          7192 => x"84",
          7193 => x"95",
          7194 => x"84",
          7195 => x"84",
          7196 => x"a0",
          7197 => x"b8",
          7198 => x"80",
          7199 => x"52",
          7200 => x"51",
          7201 => x"3f",
          7202 => x"08",
          7203 => x"34",
          7204 => x"1f",
          7205 => x"d4",
          7206 => x"84",
          7207 => x"0b",
          7208 => x"84",
          7209 => x"5c",
          7210 => x"34",
          7211 => x"1d",
          7212 => x"d4",
          7213 => x"d0",
          7214 => x"fe",
          7215 => x"70",
          7216 => x"06",
          7217 => x"5c",
          7218 => x"78",
          7219 => x"77",
          7220 => x"84",
          7221 => x"70",
          7222 => x"84",
          7223 => x"05",
          7224 => x"56",
          7225 => x"34",
          7226 => x"15",
          7227 => x"d4",
          7228 => x"fa",
          7229 => x"80",
          7230 => x"38",
          7231 => x"80",
          7232 => x"38",
          7233 => x"9b",
          7234 => x"e4",
          7235 => x"e4",
          7236 => x"0d",
          7237 => x"84",
          7238 => x"71",
          7239 => x"11",
          7240 => x"05",
          7241 => x"12",
          7242 => x"2b",
          7243 => x"ff",
          7244 => x"2a",
          7245 => x"5e",
          7246 => x"34",
          7247 => x"34",
          7248 => x"d4",
          7249 => x"88",
          7250 => x"75",
          7251 => x"7b",
          7252 => x"84",
          7253 => x"70",
          7254 => x"81",
          7255 => x"88",
          7256 => x"83",
          7257 => x"f8",
          7258 => x"64",
          7259 => x"06",
          7260 => x"4a",
          7261 => x"5e",
          7262 => x"63",
          7263 => x"76",
          7264 => x"41",
          7265 => x"05",
          7266 => x"d4",
          7267 => x"63",
          7268 => x"81",
          7269 => x"84",
          7270 => x"05",
          7271 => x"ed",
          7272 => x"54",
          7273 => x"7b",
          7274 => x"83",
          7275 => x"42",
          7276 => x"39",
          7277 => x"ff",
          7278 => x"70",
          7279 => x"06",
          7280 => x"83",
          7281 => x"88",
          7282 => x"10",
          7283 => x"70",
          7284 => x"33",
          7285 => x"71",
          7286 => x"53",
          7287 => x"58",
          7288 => x"73",
          7289 => x"f7",
          7290 => x"39",
          7291 => x"fa",
          7292 => x"7a",
          7293 => x"38",
          7294 => x"ff",
          7295 => x"7b",
          7296 => x"38",
          7297 => x"84",
          7298 => x"84",
          7299 => x"a0",
          7300 => x"b8",
          7301 => x"80",
          7302 => x"52",
          7303 => x"51",
          7304 => x"3f",
          7305 => x"08",
          7306 => x"34",
          7307 => x"1b",
          7308 => x"d4",
          7309 => x"84",
          7310 => x"0b",
          7311 => x"84",
          7312 => x"58",
          7313 => x"34",
          7314 => x"19",
          7315 => x"d4",
          7316 => x"d0",
          7317 => x"fe",
          7318 => x"70",
          7319 => x"06",
          7320 => x"58",
          7321 => x"74",
          7322 => x"34",
          7323 => x"05",
          7324 => x"d0",
          7325 => x"10",
          7326 => x"d4",
          7327 => x"05",
          7328 => x"61",
          7329 => x"81",
          7330 => x"34",
          7331 => x"80",
          7332 => x"de",
          7333 => x"ff",
          7334 => x"61",
          7335 => x"c0",
          7336 => x"39",
          7337 => x"82",
          7338 => x"51",
          7339 => x"7f",
          7340 => x"b8",
          7341 => x"3d",
          7342 => x"1e",
          7343 => x"83",
          7344 => x"8b",
          7345 => x"2b",
          7346 => x"86",
          7347 => x"12",
          7348 => x"2b",
          7349 => x"07",
          7350 => x"14",
          7351 => x"33",
          7352 => x"07",
          7353 => x"43",
          7354 => x"5b",
          7355 => x"5c",
          7356 => x"64",
          7357 => x"7a",
          7358 => x"34",
          7359 => x"08",
          7360 => x"11",
          7361 => x"33",
          7362 => x"71",
          7363 => x"74",
          7364 => x"33",
          7365 => x"71",
          7366 => x"70",
          7367 => x"41",
          7368 => x"59",
          7369 => x"64",
          7370 => x"7a",
          7371 => x"34",
          7372 => x"08",
          7373 => x"81",
          7374 => x"88",
          7375 => x"ff",
          7376 => x"88",
          7377 => x"5a",
          7378 => x"34",
          7379 => x"34",
          7380 => x"08",
          7381 => x"11",
          7382 => x"33",
          7383 => x"71",
          7384 => x"74",
          7385 => x"81",
          7386 => x"88",
          7387 => x"88",
          7388 => x"5e",
          7389 => x"45",
          7390 => x"34",
          7391 => x"34",
          7392 => x"08",
          7393 => x"33",
          7394 => x"71",
          7395 => x"83",
          7396 => x"05",
          7397 => x"83",
          7398 => x"88",
          7399 => x"88",
          7400 => x"40",
          7401 => x"55",
          7402 => x"18",
          7403 => x"18",
          7404 => x"d4",
          7405 => x"82",
          7406 => x"12",
          7407 => x"2b",
          7408 => x"62",
          7409 => x"2b",
          7410 => x"5d",
          7411 => x"05",
          7412 => x"ef",
          7413 => x"d4",
          7414 => x"05",
          7415 => x"ff",
          7416 => x"fc",
          7417 => x"ff",
          7418 => x"b8",
          7419 => x"80",
          7420 => x"d0",
          7421 => x"80",
          7422 => x"84",
          7423 => x"fe",
          7424 => x"84",
          7425 => x"56",
          7426 => x"81",
          7427 => x"34",
          7428 => x"08",
          7429 => x"16",
          7430 => x"85",
          7431 => x"b8",
          7432 => x"7f",
          7433 => x"81",
          7434 => x"34",
          7435 => x"08",
          7436 => x"22",
          7437 => x"80",
          7438 => x"83",
          7439 => x"70",
          7440 => x"43",
          7441 => x"88",
          7442 => x"89",
          7443 => x"b8",
          7444 => x"10",
          7445 => x"b8",
          7446 => x"f8",
          7447 => x"7f",
          7448 => x"81",
          7449 => x"34",
          7450 => x"bd",
          7451 => x"fc",
          7452 => x"19",
          7453 => x"33",
          7454 => x"71",
          7455 => x"79",
          7456 => x"33",
          7457 => x"71",
          7458 => x"70",
          7459 => x"48",
          7460 => x"55",
          7461 => x"05",
          7462 => x"85",
          7463 => x"b8",
          7464 => x"1e",
          7465 => x"85",
          7466 => x"8b",
          7467 => x"2b",
          7468 => x"86",
          7469 => x"15",
          7470 => x"2b",
          7471 => x"2a",
          7472 => x"48",
          7473 => x"40",
          7474 => x"05",
          7475 => x"87",
          7476 => x"b8",
          7477 => x"70",
          7478 => x"33",
          7479 => x"07",
          7480 => x"06",
          7481 => x"59",
          7482 => x"75",
          7483 => x"81",
          7484 => x"b8",
          7485 => x"1f",
          7486 => x"12",
          7487 => x"2b",
          7488 => x"07",
          7489 => x"33",
          7490 => x"71",
          7491 => x"70",
          7492 => x"ff",
          7493 => x"05",
          7494 => x"48",
          7495 => x"5d",
          7496 => x"41",
          7497 => x"34",
          7498 => x"34",
          7499 => x"08",
          7500 => x"33",
          7501 => x"71",
          7502 => x"83",
          7503 => x"05",
          7504 => x"12",
          7505 => x"2b",
          7506 => x"ff",
          7507 => x"2a",
          7508 => x"5e",
          7509 => x"5b",
          7510 => x"76",
          7511 => x"34",
          7512 => x"ff",
          7513 => x"b3",
          7514 => x"33",
          7515 => x"71",
          7516 => x"83",
          7517 => x"05",
          7518 => x"85",
          7519 => x"88",
          7520 => x"88",
          7521 => x"5a",
          7522 => x"78",
          7523 => x"79",
          7524 => x"84",
          7525 => x"70",
          7526 => x"33",
          7527 => x"71",
          7528 => x"83",
          7529 => x"05",
          7530 => x"87",
          7531 => x"88",
          7532 => x"88",
          7533 => x"5e",
          7534 => x"55",
          7535 => x"86",
          7536 => x"60",
          7537 => x"84",
          7538 => x"18",
          7539 => x"12",
          7540 => x"2b",
          7541 => x"ff",
          7542 => x"2a",
          7543 => x"55",
          7544 => x"78",
          7545 => x"84",
          7546 => x"70",
          7547 => x"81",
          7548 => x"8b",
          7549 => x"2b",
          7550 => x"70",
          7551 => x"33",
          7552 => x"07",
          7553 => x"8f",
          7554 => x"77",
          7555 => x"2a",
          7556 => x"5f",
          7557 => x"5e",
          7558 => x"17",
          7559 => x"17",
          7560 => x"d4",
          7561 => x"70",
          7562 => x"33",
          7563 => x"71",
          7564 => x"74",
          7565 => x"81",
          7566 => x"88",
          7567 => x"ff",
          7568 => x"88",
          7569 => x"5e",
          7570 => x"5d",
          7571 => x"34",
          7572 => x"34",
          7573 => x"08",
          7574 => x"11",
          7575 => x"33",
          7576 => x"71",
          7577 => x"74",
          7578 => x"33",
          7579 => x"71",
          7580 => x"83",
          7581 => x"05",
          7582 => x"85",
          7583 => x"88",
          7584 => x"88",
          7585 => x"49",
          7586 => x"59",
          7587 => x"57",
          7588 => x"1d",
          7589 => x"1d",
          7590 => x"d4",
          7591 => x"84",
          7592 => x"12",
          7593 => x"2b",
          7594 => x"07",
          7595 => x"14",
          7596 => x"33",
          7597 => x"07",
          7598 => x"5f",
          7599 => x"40",
          7600 => x"77",
          7601 => x"7b",
          7602 => x"84",
          7603 => x"16",
          7604 => x"12",
          7605 => x"2b",
          7606 => x"ff",
          7607 => x"2a",
          7608 => x"59",
          7609 => x"79",
          7610 => x"84",
          7611 => x"70",
          7612 => x"33",
          7613 => x"71",
          7614 => x"83",
          7615 => x"05",
          7616 => x"15",
          7617 => x"2b",
          7618 => x"2a",
          7619 => x"5d",
          7620 => x"55",
          7621 => x"75",
          7622 => x"84",
          7623 => x"70",
          7624 => x"81",
          7625 => x"8b",
          7626 => x"2b",
          7627 => x"82",
          7628 => x"15",
          7629 => x"2b",
          7630 => x"2a",
          7631 => x"5d",
          7632 => x"55",
          7633 => x"34",
          7634 => x"34",
          7635 => x"08",
          7636 => x"11",
          7637 => x"33",
          7638 => x"07",
          7639 => x"56",
          7640 => x"42",
          7641 => x"7e",
          7642 => x"51",
          7643 => x"3f",
          7644 => x"08",
          7645 => x"61",
          7646 => x"70",
          7647 => x"06",
          7648 => x"f1",
          7649 => x"19",
          7650 => x"33",
          7651 => x"71",
          7652 => x"79",
          7653 => x"33",
          7654 => x"71",
          7655 => x"70",
          7656 => x"48",
          7657 => x"55",
          7658 => x"05",
          7659 => x"85",
          7660 => x"b8",
          7661 => x"1e",
          7662 => x"85",
          7663 => x"8b",
          7664 => x"2b",
          7665 => x"86",
          7666 => x"15",
          7667 => x"2b",
          7668 => x"2a",
          7669 => x"48",
          7670 => x"56",
          7671 => x"05",
          7672 => x"87",
          7673 => x"b8",
          7674 => x"70",
          7675 => x"33",
          7676 => x"07",
          7677 => x"06",
          7678 => x"5c",
          7679 => x"78",
          7680 => x"81",
          7681 => x"b8",
          7682 => x"1f",
          7683 => x"12",
          7684 => x"2b",
          7685 => x"07",
          7686 => x"33",
          7687 => x"71",
          7688 => x"70",
          7689 => x"ff",
          7690 => x"05",
          7691 => x"5d",
          7692 => x"58",
          7693 => x"40",
          7694 => x"34",
          7695 => x"34",
          7696 => x"08",
          7697 => x"33",
          7698 => x"71",
          7699 => x"83",
          7700 => x"05",
          7701 => x"12",
          7702 => x"2b",
          7703 => x"ff",
          7704 => x"2a",
          7705 => x"58",
          7706 => x"5b",
          7707 => x"78",
          7708 => x"77",
          7709 => x"06",
          7710 => x"39",
          7711 => x"54",
          7712 => x"84",
          7713 => x"5f",
          7714 => x"08",
          7715 => x"38",
          7716 => x"52",
          7717 => x"08",
          7718 => x"cf",
          7719 => x"df",
          7720 => x"5b",
          7721 => x"ef",
          7722 => x"e9",
          7723 => x"0d",
          7724 => x"84",
          7725 => x"58",
          7726 => x"2e",
          7727 => x"54",
          7728 => x"73",
          7729 => x"0c",
          7730 => x"04",
          7731 => x"d3",
          7732 => x"e4",
          7733 => x"b8",
          7734 => x"2e",
          7735 => x"53",
          7736 => x"b8",
          7737 => x"fe",
          7738 => x"73",
          7739 => x"0c",
          7740 => x"04",
          7741 => x"0b",
          7742 => x"0c",
          7743 => x"84",
          7744 => x"82",
          7745 => x"76",
          7746 => x"f4",
          7747 => x"f0",
          7748 => x"d4",
          7749 => x"75",
          7750 => x"81",
          7751 => x"b8",
          7752 => x"76",
          7753 => x"81",
          7754 => x"34",
          7755 => x"08",
          7756 => x"17",
          7757 => x"87",
          7758 => x"b8",
          7759 => x"b8",
          7760 => x"05",
          7761 => x"07",
          7762 => x"ff",
          7763 => x"2a",
          7764 => x"56",
          7765 => x"34",
          7766 => x"34",
          7767 => x"22",
          7768 => x"10",
          7769 => x"08",
          7770 => x"55",
          7771 => x"15",
          7772 => x"83",
          7773 => x"54",
          7774 => x"fe",
          7775 => x"cc",
          7776 => x"0d",
          7777 => x"33",
          7778 => x"70",
          7779 => x"38",
          7780 => x"11",
          7781 => x"84",
          7782 => x"83",
          7783 => x"fe",
          7784 => x"93",
          7785 => x"83",
          7786 => x"26",
          7787 => x"51",
          7788 => x"84",
          7789 => x"81",
          7790 => x"72",
          7791 => x"84",
          7792 => x"34",
          7793 => x"12",
          7794 => x"84",
          7795 => x"84",
          7796 => x"f7",
          7797 => x"7e",
          7798 => x"05",
          7799 => x"5a",
          7800 => x"81",
          7801 => x"26",
          7802 => x"b8",
          7803 => x"54",
          7804 => x"54",
          7805 => x"bd",
          7806 => x"85",
          7807 => x"98",
          7808 => x"53",
          7809 => x"51",
          7810 => x"84",
          7811 => x"81",
          7812 => x"74",
          7813 => x"38",
          7814 => x"8c",
          7815 => x"e2",
          7816 => x"26",
          7817 => x"fc",
          7818 => x"54",
          7819 => x"83",
          7820 => x"73",
          7821 => x"b8",
          7822 => x"3d",
          7823 => x"80",
          7824 => x"70",
          7825 => x"5a",
          7826 => x"78",
          7827 => x"38",
          7828 => x"3d",
          7829 => x"60",
          7830 => x"af",
          7831 => x"5c",
          7832 => x"54",
          7833 => x"87",
          7834 => x"e0",
          7835 => x"73",
          7836 => x"83",
          7837 => x"38",
          7838 => x"0b",
          7839 => x"8c",
          7840 => x"75",
          7841 => x"d7",
          7842 => x"b8",
          7843 => x"ff",
          7844 => x"80",
          7845 => x"87",
          7846 => x"08",
          7847 => x"38",
          7848 => x"d6",
          7849 => x"80",
          7850 => x"73",
          7851 => x"38",
          7852 => x"55",
          7853 => x"e4",
          7854 => x"0d",
          7855 => x"16",
          7856 => x"81",
          7857 => x"55",
          7858 => x"26",
          7859 => x"d5",
          7860 => x"0d",
          7861 => x"05",
          7862 => x"02",
          7863 => x"05",
          7864 => x"55",
          7865 => x"73",
          7866 => x"84",
          7867 => x"33",
          7868 => x"06",
          7869 => x"73",
          7870 => x"0b",
          7871 => x"8c",
          7872 => x"70",
          7873 => x"38",
          7874 => x"ad",
          7875 => x"2e",
          7876 => x"53",
          7877 => x"e4",
          7878 => x"0d",
          7879 => x"0a",
          7880 => x"84",
          7881 => x"86",
          7882 => x"81",
          7883 => x"80",
          7884 => x"e4",
          7885 => x"0d",
          7886 => x"2b",
          7887 => x"8c",
          7888 => x"70",
          7889 => x"08",
          7890 => x"81",
          7891 => x"70",
          7892 => x"38",
          7893 => x"8c",
          7894 => x"ea",
          7895 => x"98",
          7896 => x"70",
          7897 => x"72",
          7898 => x"92",
          7899 => x"71",
          7900 => x"54",
          7901 => x"ff",
          7902 => x"08",
          7903 => x"73",
          7904 => x"90",
          7905 => x"0d",
          7906 => x"0b",
          7907 => x"71",
          7908 => x"74",
          7909 => x"81",
          7910 => x"77",
          7911 => x"83",
          7912 => x"38",
          7913 => x"52",
          7914 => x"51",
          7915 => x"84",
          7916 => x"80",
          7917 => x"81",
          7918 => x"b8",
          7919 => x"3d",
          7920 => x"54",
          7921 => x"53",
          7922 => x"53",
          7923 => x"52",
          7924 => x"3f",
          7925 => x"b8",
          7926 => x"2e",
          7927 => x"d9",
          7928 => x"e4",
          7929 => x"34",
          7930 => x"70",
          7931 => x"31",
          7932 => x"84",
          7933 => x"5c",
          7934 => x"74",
          7935 => x"9b",
          7936 => x"33",
          7937 => x"2e",
          7938 => x"ff",
          7939 => x"54",
          7940 => x"79",
          7941 => x"33",
          7942 => x"3f",
          7943 => x"57",
          7944 => x"2e",
          7945 => x"fe",
          7946 => x"18",
          7947 => x"81",
          7948 => x"06",
          7949 => x"b8",
          7950 => x"80",
          7951 => x"80",
          7952 => x"05",
          7953 => x"17",
          7954 => x"38",
          7955 => x"84",
          7956 => x"ff",
          7957 => x"b7",
          7958 => x"d2",
          7959 => x"d2",
          7960 => x"34",
          7961 => x"ba",
          7962 => x"c1",
          7963 => x"34",
          7964 => x"84",
          7965 => x"80",
          7966 => x"9d",
          7967 => x"c1",
          7968 => x"19",
          7969 => x"0b",
          7970 => x"34",
          7971 => x"55",
          7972 => x"19",
          7973 => x"2a",
          7974 => x"a1",
          7975 => x"90",
          7976 => x"84",
          7977 => x"74",
          7978 => x"7a",
          7979 => x"34",
          7980 => x"5b",
          7981 => x"19",
          7982 => x"2a",
          7983 => x"a5",
          7984 => x"90",
          7985 => x"84",
          7986 => x"7a",
          7987 => x"74",
          7988 => x"34",
          7989 => x"81",
          7990 => x"1a",
          7991 => x"54",
          7992 => x"52",
          7993 => x"51",
          7994 => x"76",
          7995 => x"80",
          7996 => x"81",
          7997 => x"fb",
          7998 => x"b8",
          7999 => x"2e",
          8000 => x"fd",
          8001 => x"3d",
          8002 => x"70",
          8003 => x"56",
          8004 => x"88",
          8005 => x"08",
          8006 => x"38",
          8007 => x"84",
          8008 => x"8f",
          8009 => x"ff",
          8010 => x"58",
          8011 => x"81",
          8012 => x"82",
          8013 => x"38",
          8014 => x"09",
          8015 => x"38",
          8016 => x"16",
          8017 => x"a8",
          8018 => x"5a",
          8019 => x"b4",
          8020 => x"2e",
          8021 => x"17",
          8022 => x"7b",
          8023 => x"06",
          8024 => x"81",
          8025 => x"b8",
          8026 => x"17",
          8027 => x"e3",
          8028 => x"e4",
          8029 => x"85",
          8030 => x"81",
          8031 => x"18",
          8032 => x"9a",
          8033 => x"ff",
          8034 => x"11",
          8035 => x"70",
          8036 => x"1b",
          8037 => x"5d",
          8038 => x"17",
          8039 => x"b5",
          8040 => x"83",
          8041 => x"5c",
          8042 => x"7d",
          8043 => x"06",
          8044 => x"81",
          8045 => x"b8",
          8046 => x"17",
          8047 => x"93",
          8048 => x"e4",
          8049 => x"85",
          8050 => x"81",
          8051 => x"18",
          8052 => x"ca",
          8053 => x"ff",
          8054 => x"11",
          8055 => x"2b",
          8056 => x"81",
          8057 => x"2a",
          8058 => x"59",
          8059 => x"ae",
          8060 => x"ff",
          8061 => x"e4",
          8062 => x"0d",
          8063 => x"2a",
          8064 => x"05",
          8065 => x"08",
          8066 => x"38",
          8067 => x"18",
          8068 => x"5d",
          8069 => x"2e",
          8070 => x"81",
          8071 => x"54",
          8072 => x"17",
          8073 => x"33",
          8074 => x"3f",
          8075 => x"08",
          8076 => x"38",
          8077 => x"5a",
          8078 => x"0c",
          8079 => x"38",
          8080 => x"fe",
          8081 => x"b8",
          8082 => x"33",
          8083 => x"88",
          8084 => x"b8",
          8085 => x"5b",
          8086 => x"04",
          8087 => x"09",
          8088 => x"b8",
          8089 => x"2a",
          8090 => x"05",
          8091 => x"08",
          8092 => x"38",
          8093 => x"18",
          8094 => x"5e",
          8095 => x"2e",
          8096 => x"82",
          8097 => x"54",
          8098 => x"17",
          8099 => x"33",
          8100 => x"3f",
          8101 => x"08",
          8102 => x"38",
          8103 => x"5a",
          8104 => x"0c",
          8105 => x"38",
          8106 => x"83",
          8107 => x"05",
          8108 => x"11",
          8109 => x"33",
          8110 => x"71",
          8111 => x"81",
          8112 => x"72",
          8113 => x"75",
          8114 => x"ff",
          8115 => x"06",
          8116 => x"e4",
          8117 => x"5e",
          8118 => x"8f",
          8119 => x"81",
          8120 => x"08",
          8121 => x"70",
          8122 => x"33",
          8123 => x"e2",
          8124 => x"84",
          8125 => x"7b",
          8126 => x"06",
          8127 => x"84",
          8128 => x"83",
          8129 => x"17",
          8130 => x"08",
          8131 => x"e4",
          8132 => x"7d",
          8133 => x"27",
          8134 => x"82",
          8135 => x"74",
          8136 => x"81",
          8137 => x"38",
          8138 => x"17",
          8139 => x"08",
          8140 => x"52",
          8141 => x"51",
          8142 => x"7a",
          8143 => x"39",
          8144 => x"17",
          8145 => x"17",
          8146 => x"18",
          8147 => x"f6",
          8148 => x"b8",
          8149 => x"2e",
          8150 => x"82",
          8151 => x"b8",
          8152 => x"18",
          8153 => x"08",
          8154 => x"31",
          8155 => x"18",
          8156 => x"38",
          8157 => x"5e",
          8158 => x"81",
          8159 => x"b8",
          8160 => x"fb",
          8161 => x"54",
          8162 => x"53",
          8163 => x"53",
          8164 => x"52",
          8165 => x"3f",
          8166 => x"b8",
          8167 => x"2e",
          8168 => x"fd",
          8169 => x"b8",
          8170 => x"18",
          8171 => x"08",
          8172 => x"31",
          8173 => x"08",
          8174 => x"a0",
          8175 => x"fd",
          8176 => x"17",
          8177 => x"82",
          8178 => x"06",
          8179 => x"81",
          8180 => x"08",
          8181 => x"05",
          8182 => x"81",
          8183 => x"f4",
          8184 => x"5a",
          8185 => x"81",
          8186 => x"08",
          8187 => x"70",
          8188 => x"33",
          8189 => x"da",
          8190 => x"84",
          8191 => x"7d",
          8192 => x"06",
          8193 => x"84",
          8194 => x"83",
          8195 => x"17",
          8196 => x"08",
          8197 => x"e4",
          8198 => x"74",
          8199 => x"27",
          8200 => x"82",
          8201 => x"74",
          8202 => x"81",
          8203 => x"38",
          8204 => x"17",
          8205 => x"08",
          8206 => x"52",
          8207 => x"51",
          8208 => x"7c",
          8209 => x"39",
          8210 => x"17",
          8211 => x"08",
          8212 => x"52",
          8213 => x"51",
          8214 => x"fa",
          8215 => x"5b",
          8216 => x"38",
          8217 => x"f2",
          8218 => x"62",
          8219 => x"59",
          8220 => x"76",
          8221 => x"75",
          8222 => x"27",
          8223 => x"33",
          8224 => x"2e",
          8225 => x"78",
          8226 => x"38",
          8227 => x"82",
          8228 => x"84",
          8229 => x"90",
          8230 => x"75",
          8231 => x"1a",
          8232 => x"80",
          8233 => x"08",
          8234 => x"78",
          8235 => x"38",
          8236 => x"7c",
          8237 => x"7c",
          8238 => x"06",
          8239 => x"81",
          8240 => x"b8",
          8241 => x"19",
          8242 => x"87",
          8243 => x"e4",
          8244 => x"85",
          8245 => x"81",
          8246 => x"1a",
          8247 => x"79",
          8248 => x"75",
          8249 => x"06",
          8250 => x"83",
          8251 => x"58",
          8252 => x"1f",
          8253 => x"2a",
          8254 => x"1f",
          8255 => x"83",
          8256 => x"84",
          8257 => x"90",
          8258 => x"74",
          8259 => x"81",
          8260 => x"38",
          8261 => x"a8",
          8262 => x"58",
          8263 => x"1a",
          8264 => x"76",
          8265 => x"e1",
          8266 => x"33",
          8267 => x"7c",
          8268 => x"81",
          8269 => x"38",
          8270 => x"53",
          8271 => x"81",
          8272 => x"f1",
          8273 => x"b8",
          8274 => x"2e",
          8275 => x"58",
          8276 => x"b4",
          8277 => x"58",
          8278 => x"38",
          8279 => x"83",
          8280 => x"05",
          8281 => x"11",
          8282 => x"2b",
          8283 => x"7e",
          8284 => x"07",
          8285 => x"5c",
          8286 => x"7d",
          8287 => x"75",
          8288 => x"7d",
          8289 => x"79",
          8290 => x"7d",
          8291 => x"7a",
          8292 => x"81",
          8293 => x"34",
          8294 => x"75",
          8295 => x"70",
          8296 => x"1b",
          8297 => x"1b",
          8298 => x"5a",
          8299 => x"b7",
          8300 => x"83",
          8301 => x"5e",
          8302 => x"7d",
          8303 => x"06",
          8304 => x"81",
          8305 => x"b8",
          8306 => x"19",
          8307 => x"83",
          8308 => x"e4",
          8309 => x"85",
          8310 => x"81",
          8311 => x"1a",
          8312 => x"7b",
          8313 => x"79",
          8314 => x"19",
          8315 => x"1b",
          8316 => x"5f",
          8317 => x"55",
          8318 => x"8f",
          8319 => x"2b",
          8320 => x"77",
          8321 => x"71",
          8322 => x"74",
          8323 => x"0b",
          8324 => x"7d",
          8325 => x"1a",
          8326 => x"80",
          8327 => x"08",
          8328 => x"76",
          8329 => x"38",
          8330 => x"53",
          8331 => x"53",
          8332 => x"52",
          8333 => x"3f",
          8334 => x"b8",
          8335 => x"2e",
          8336 => x"80",
          8337 => x"b8",
          8338 => x"1a",
          8339 => x"08",
          8340 => x"08",
          8341 => x"08",
          8342 => x"08",
          8343 => x"5c",
          8344 => x"8b",
          8345 => x"33",
          8346 => x"2e",
          8347 => x"81",
          8348 => x"76",
          8349 => x"33",
          8350 => x"3f",
          8351 => x"08",
          8352 => x"38",
          8353 => x"58",
          8354 => x"0c",
          8355 => x"38",
          8356 => x"06",
          8357 => x"7b",
          8358 => x"56",
          8359 => x"7a",
          8360 => x"33",
          8361 => x"71",
          8362 => x"56",
          8363 => x"34",
          8364 => x"1a",
          8365 => x"39",
          8366 => x"53",
          8367 => x"53",
          8368 => x"52",
          8369 => x"3f",
          8370 => x"b8",
          8371 => x"2e",
          8372 => x"fc",
          8373 => x"b8",
          8374 => x"1a",
          8375 => x"08",
          8376 => x"08",
          8377 => x"08",
          8378 => x"08",
          8379 => x"5e",
          8380 => x"fb",
          8381 => x"19",
          8382 => x"82",
          8383 => x"06",
          8384 => x"81",
          8385 => x"53",
          8386 => x"19",
          8387 => x"c2",
          8388 => x"fb",
          8389 => x"54",
          8390 => x"19",
          8391 => x"1a",
          8392 => x"ee",
          8393 => x"5c",
          8394 => x"08",
          8395 => x"81",
          8396 => x"38",
          8397 => x"08",
          8398 => x"b4",
          8399 => x"a8",
          8400 => x"a0",
          8401 => x"b8",
          8402 => x"40",
          8403 => x"7e",
          8404 => x"38",
          8405 => x"55",
          8406 => x"09",
          8407 => x"e3",
          8408 => x"7d",
          8409 => x"52",
          8410 => x"51",
          8411 => x"7c",
          8412 => x"39",
          8413 => x"53",
          8414 => x"53",
          8415 => x"52",
          8416 => x"3f",
          8417 => x"b8",
          8418 => x"2e",
          8419 => x"fb",
          8420 => x"b8",
          8421 => x"1a",
          8422 => x"08",
          8423 => x"08",
          8424 => x"08",
          8425 => x"08",
          8426 => x"5e",
          8427 => x"fb",
          8428 => x"19",
          8429 => x"82",
          8430 => x"06",
          8431 => x"81",
          8432 => x"53",
          8433 => x"19",
          8434 => x"86",
          8435 => x"fa",
          8436 => x"54",
          8437 => x"76",
          8438 => x"33",
          8439 => x"3f",
          8440 => x"8b",
          8441 => x"10",
          8442 => x"7a",
          8443 => x"ff",
          8444 => x"5f",
          8445 => x"1f",
          8446 => x"2a",
          8447 => x"1f",
          8448 => x"39",
          8449 => x"88",
          8450 => x"82",
          8451 => x"06",
          8452 => x"11",
          8453 => x"70",
          8454 => x"0a",
          8455 => x"0a",
          8456 => x"58",
          8457 => x"7d",
          8458 => x"88",
          8459 => x"b9",
          8460 => x"90",
          8461 => x"ba",
          8462 => x"98",
          8463 => x"bb",
          8464 => x"cf",
          8465 => x"0d",
          8466 => x"08",
          8467 => x"7a",
          8468 => x"90",
          8469 => x"76",
          8470 => x"f4",
          8471 => x"1a",
          8472 => x"ec",
          8473 => x"08",
          8474 => x"73",
          8475 => x"d7",
          8476 => x"2e",
          8477 => x"76",
          8478 => x"56",
          8479 => x"76",
          8480 => x"82",
          8481 => x"26",
          8482 => x"75",
          8483 => x"f0",
          8484 => x"b8",
          8485 => x"2e",
          8486 => x"80",
          8487 => x"e4",
          8488 => x"b1",
          8489 => x"e4",
          8490 => x"30",
          8491 => x"80",
          8492 => x"07",
          8493 => x"55",
          8494 => x"38",
          8495 => x"09",
          8496 => x"b5",
          8497 => x"74",
          8498 => x"0c",
          8499 => x"04",
          8500 => x"91",
          8501 => x"e4",
          8502 => x"39",
          8503 => x"51",
          8504 => x"81",
          8505 => x"b8",
          8506 => x"db",
          8507 => x"e4",
          8508 => x"b8",
          8509 => x"2e",
          8510 => x"19",
          8511 => x"e4",
          8512 => x"38",
          8513 => x"dd",
          8514 => x"56",
          8515 => x"76",
          8516 => x"82",
          8517 => x"79",
          8518 => x"3f",
          8519 => x"b8",
          8520 => x"2e",
          8521 => x"84",
          8522 => x"09",
          8523 => x"72",
          8524 => x"70",
          8525 => x"b8",
          8526 => x"51",
          8527 => x"73",
          8528 => x"84",
          8529 => x"80",
          8530 => x"90",
          8531 => x"81",
          8532 => x"a3",
          8533 => x"1a",
          8534 => x"9b",
          8535 => x"57",
          8536 => x"39",
          8537 => x"fe",
          8538 => x"53",
          8539 => x"51",
          8540 => x"84",
          8541 => x"84",
          8542 => x"30",
          8543 => x"e4",
          8544 => x"25",
          8545 => x"7a",
          8546 => x"74",
          8547 => x"75",
          8548 => x"9c",
          8549 => x"05",
          8550 => x"56",
          8551 => x"26",
          8552 => x"15",
          8553 => x"84",
          8554 => x"07",
          8555 => x"1a",
          8556 => x"74",
          8557 => x"0c",
          8558 => x"04",
          8559 => x"b8",
          8560 => x"3d",
          8561 => x"b8",
          8562 => x"fe",
          8563 => x"80",
          8564 => x"38",
          8565 => x"52",
          8566 => x"8b",
          8567 => x"e4",
          8568 => x"a7",
          8569 => x"e4",
          8570 => x"e4",
          8571 => x"0d",
          8572 => x"74",
          8573 => x"b9",
          8574 => x"ff",
          8575 => x"3d",
          8576 => x"71",
          8577 => x"58",
          8578 => x"0a",
          8579 => x"38",
          8580 => x"53",
          8581 => x"38",
          8582 => x"0c",
          8583 => x"55",
          8584 => x"38",
          8585 => x"75",
          8586 => x"cc",
          8587 => x"2a",
          8588 => x"88",
          8589 => x"56",
          8590 => x"a9",
          8591 => x"08",
          8592 => x"74",
          8593 => x"98",
          8594 => x"82",
          8595 => x"2e",
          8596 => x"89",
          8597 => x"19",
          8598 => x"ff",
          8599 => x"05",
          8600 => x"80",
          8601 => x"b8",
          8602 => x"3d",
          8603 => x"0b",
          8604 => x"0c",
          8605 => x"04",
          8606 => x"55",
          8607 => x"ff",
          8608 => x"17",
          8609 => x"2b",
          8610 => x"76",
          8611 => x"9c",
          8612 => x"fe",
          8613 => x"54",
          8614 => x"75",
          8615 => x"38",
          8616 => x"76",
          8617 => x"19",
          8618 => x"53",
          8619 => x"0c",
          8620 => x"74",
          8621 => x"ec",
          8622 => x"b8",
          8623 => x"84",
          8624 => x"ff",
          8625 => x"81",
          8626 => x"e4",
          8627 => x"9e",
          8628 => x"08",
          8629 => x"e4",
          8630 => x"ff",
          8631 => x"76",
          8632 => x"76",
          8633 => x"ff",
          8634 => x"0b",
          8635 => x"0c",
          8636 => x"04",
          8637 => x"7f",
          8638 => x"12",
          8639 => x"5c",
          8640 => x"80",
          8641 => x"86",
          8642 => x"98",
          8643 => x"17",
          8644 => x"56",
          8645 => x"b2",
          8646 => x"ff",
          8647 => x"9d",
          8648 => x"94",
          8649 => x"58",
          8650 => x"79",
          8651 => x"1a",
          8652 => x"74",
          8653 => x"f5",
          8654 => x"18",
          8655 => x"18",
          8656 => x"b8",
          8657 => x"0c",
          8658 => x"84",
          8659 => x"8f",
          8660 => x"77",
          8661 => x"8a",
          8662 => x"05",
          8663 => x"06",
          8664 => x"38",
          8665 => x"51",
          8666 => x"84",
          8667 => x"5d",
          8668 => x"0b",
          8669 => x"08",
          8670 => x"81",
          8671 => x"e4",
          8672 => x"c6",
          8673 => x"08",
          8674 => x"08",
          8675 => x"38",
          8676 => x"81",
          8677 => x"17",
          8678 => x"51",
          8679 => x"84",
          8680 => x"5d",
          8681 => x"b8",
          8682 => x"2e",
          8683 => x"82",
          8684 => x"e4",
          8685 => x"ff",
          8686 => x"56",
          8687 => x"08",
          8688 => x"86",
          8689 => x"e4",
          8690 => x"33",
          8691 => x"80",
          8692 => x"18",
          8693 => x"fe",
          8694 => x"80",
          8695 => x"27",
          8696 => x"19",
          8697 => x"29",
          8698 => x"05",
          8699 => x"b4",
          8700 => x"19",
          8701 => x"78",
          8702 => x"76",
          8703 => x"58",
          8704 => x"55",
          8705 => x"74",
          8706 => x"22",
          8707 => x"27",
          8708 => x"81",
          8709 => x"53",
          8710 => x"19",
          8711 => x"b2",
          8712 => x"e4",
          8713 => x"38",
          8714 => x"dd",
          8715 => x"18",
          8716 => x"84",
          8717 => x"8f",
          8718 => x"75",
          8719 => x"08",
          8720 => x"70",
          8721 => x"33",
          8722 => x"86",
          8723 => x"e4",
          8724 => x"38",
          8725 => x"08",
          8726 => x"b4",
          8727 => x"1a",
          8728 => x"74",
          8729 => x"27",
          8730 => x"82",
          8731 => x"7b",
          8732 => x"81",
          8733 => x"38",
          8734 => x"19",
          8735 => x"08",
          8736 => x"52",
          8737 => x"51",
          8738 => x"fe",
          8739 => x"19",
          8740 => x"83",
          8741 => x"55",
          8742 => x"09",
          8743 => x"38",
          8744 => x"0c",
          8745 => x"1a",
          8746 => x"5e",
          8747 => x"75",
          8748 => x"85",
          8749 => x"22",
          8750 => x"b0",
          8751 => x"98",
          8752 => x"fc",
          8753 => x"0b",
          8754 => x"0c",
          8755 => x"04",
          8756 => x"64",
          8757 => x"84",
          8758 => x"5b",
          8759 => x"98",
          8760 => x"5e",
          8761 => x"2e",
          8762 => x"b8",
          8763 => x"5a",
          8764 => x"19",
          8765 => x"82",
          8766 => x"19",
          8767 => x"55",
          8768 => x"09",
          8769 => x"94",
          8770 => x"75",
          8771 => x"52",
          8772 => x"51",
          8773 => x"84",
          8774 => x"80",
          8775 => x"ff",
          8776 => x"79",
          8777 => x"76",
          8778 => x"90",
          8779 => x"08",
          8780 => x"58",
          8781 => x"82",
          8782 => x"18",
          8783 => x"70",
          8784 => x"5b",
          8785 => x"1d",
          8786 => x"e5",
          8787 => x"78",
          8788 => x"30",
          8789 => x"71",
          8790 => x"54",
          8791 => x"55",
          8792 => x"74",
          8793 => x"43",
          8794 => x"2e",
          8795 => x"75",
          8796 => x"86",
          8797 => x"5d",
          8798 => x"51",
          8799 => x"84",
          8800 => x"5b",
          8801 => x"08",
          8802 => x"98",
          8803 => x"75",
          8804 => x"7a",
          8805 => x"0c",
          8806 => x"04",
          8807 => x"19",
          8808 => x"52",
          8809 => x"51",
          8810 => x"81",
          8811 => x"e4",
          8812 => x"09",
          8813 => x"ef",
          8814 => x"e4",
          8815 => x"34",
          8816 => x"a8",
          8817 => x"84",
          8818 => x"58",
          8819 => x"1a",
          8820 => x"b5",
          8821 => x"33",
          8822 => x"2e",
          8823 => x"fe",
          8824 => x"54",
          8825 => x"a0",
          8826 => x"53",
          8827 => x"19",
          8828 => x"de",
          8829 => x"fe",
          8830 => x"8f",
          8831 => x"06",
          8832 => x"76",
          8833 => x"06",
          8834 => x"2e",
          8835 => x"18",
          8836 => x"bf",
          8837 => x"1f",
          8838 => x"05",
          8839 => x"5e",
          8840 => x"ab",
          8841 => x"55",
          8842 => x"cc",
          8843 => x"75",
          8844 => x"81",
          8845 => x"38",
          8846 => x"5b",
          8847 => x"1d",
          8848 => x"b8",
          8849 => x"3d",
          8850 => x"5b",
          8851 => x"8d",
          8852 => x"7d",
          8853 => x"81",
          8854 => x"8c",
          8855 => x"19",
          8856 => x"33",
          8857 => x"07",
          8858 => x"75",
          8859 => x"77",
          8860 => x"bf",
          8861 => x"f3",
          8862 => x"81",
          8863 => x"83",
          8864 => x"33",
          8865 => x"11",
          8866 => x"71",
          8867 => x"52",
          8868 => x"80",
          8869 => x"38",
          8870 => x"26",
          8871 => x"79",
          8872 => x"76",
          8873 => x"62",
          8874 => x"5a",
          8875 => x"8c",
          8876 => x"38",
          8877 => x"86",
          8878 => x"59",
          8879 => x"2e",
          8880 => x"81",
          8881 => x"dd",
          8882 => x"61",
          8883 => x"63",
          8884 => x"70",
          8885 => x"5e",
          8886 => x"39",
          8887 => x"ff",
          8888 => x"81",
          8889 => x"c0",
          8890 => x"38",
          8891 => x"57",
          8892 => x"75",
          8893 => x"05",
          8894 => x"05",
          8895 => x"7f",
          8896 => x"ff",
          8897 => x"59",
          8898 => x"e4",
          8899 => x"2e",
          8900 => x"ff",
          8901 => x"0c",
          8902 => x"e4",
          8903 => x"0d",
          8904 => x"0d",
          8905 => x"5c",
          8906 => x"7b",
          8907 => x"3f",
          8908 => x"08",
          8909 => x"e4",
          8910 => x"38",
          8911 => x"40",
          8912 => x"ac",
          8913 => x"1b",
          8914 => x"08",
          8915 => x"b4",
          8916 => x"2e",
          8917 => x"83",
          8918 => x"58",
          8919 => x"2e",
          8920 => x"81",
          8921 => x"54",
          8922 => x"1b",
          8923 => x"33",
          8924 => x"3f",
          8925 => x"08",
          8926 => x"38",
          8927 => x"57",
          8928 => x"0c",
          8929 => x"81",
          8930 => x"1c",
          8931 => x"58",
          8932 => x"2e",
          8933 => x"8b",
          8934 => x"06",
          8935 => x"06",
          8936 => x"86",
          8937 => x"81",
          8938 => x"f2",
          8939 => x"2a",
          8940 => x"75",
          8941 => x"ef",
          8942 => x"e2",
          8943 => x"2e",
          8944 => x"7c",
          8945 => x"7d",
          8946 => x"57",
          8947 => x"75",
          8948 => x"05",
          8949 => x"05",
          8950 => x"76",
          8951 => x"ff",
          8952 => x"59",
          8953 => x"e4",
          8954 => x"2e",
          8955 => x"ab",
          8956 => x"06",
          8957 => x"38",
          8958 => x"1d",
          8959 => x"70",
          8960 => x"33",
          8961 => x"05",
          8962 => x"71",
          8963 => x"5a",
          8964 => x"76",
          8965 => x"dc",
          8966 => x"2e",
          8967 => x"ff",
          8968 => x"ac",
          8969 => x"52",
          8970 => x"c8",
          8971 => x"e4",
          8972 => x"b8",
          8973 => x"2e",
          8974 => x"79",
          8975 => x"0c",
          8976 => x"04",
          8977 => x"1b",
          8978 => x"52",
          8979 => x"51",
          8980 => x"81",
          8981 => x"e4",
          8982 => x"09",
          8983 => x"a4",
          8984 => x"e4",
          8985 => x"34",
          8986 => x"a8",
          8987 => x"84",
          8988 => x"58",
          8989 => x"1c",
          8990 => x"ea",
          8991 => x"33",
          8992 => x"2e",
          8993 => x"fd",
          8994 => x"54",
          8995 => x"a0",
          8996 => x"53",
          8997 => x"1b",
          8998 => x"b6",
          8999 => x"fd",
          9000 => x"5a",
          9001 => x"ab",
          9002 => x"86",
          9003 => x"42",
          9004 => x"f2",
          9005 => x"2a",
          9006 => x"79",
          9007 => x"38",
          9008 => x"77",
          9009 => x"70",
          9010 => x"7f",
          9011 => x"59",
          9012 => x"7d",
          9013 => x"81",
          9014 => x"5d",
          9015 => x"51",
          9016 => x"84",
          9017 => x"5a",
          9018 => x"08",
          9019 => x"d9",
          9020 => x"39",
          9021 => x"fe",
          9022 => x"ff",
          9023 => x"ac",
          9024 => x"a2",
          9025 => x"33",
          9026 => x"2e",
          9027 => x"c7",
          9028 => x"08",
          9029 => x"9a",
          9030 => x"88",
          9031 => x"42",
          9032 => x"b3",
          9033 => x"70",
          9034 => x"29",
          9035 => x"55",
          9036 => x"56",
          9037 => x"18",
          9038 => x"81",
          9039 => x"33",
          9040 => x"07",
          9041 => x"75",
          9042 => x"ed",
          9043 => x"fe",
          9044 => x"38",
          9045 => x"a1",
          9046 => x"b8",
          9047 => x"10",
          9048 => x"22",
          9049 => x"1b",
          9050 => x"a0",
          9051 => x"84",
          9052 => x"2e",
          9053 => x"fe",
          9054 => x"56",
          9055 => x"8c",
          9056 => x"b0",
          9057 => x"70",
          9058 => x"06",
          9059 => x"80",
          9060 => x"74",
          9061 => x"38",
          9062 => x"05",
          9063 => x"41",
          9064 => x"38",
          9065 => x"81",
          9066 => x"5a",
          9067 => x"84",
          9068 => x"e4",
          9069 => x"0d",
          9070 => x"ff",
          9071 => x"bc",
          9072 => x"55",
          9073 => x"ea",
          9074 => x"70",
          9075 => x"13",
          9076 => x"06",
          9077 => x"5e",
          9078 => x"85",
          9079 => x"8c",
          9080 => x"22",
          9081 => x"74",
          9082 => x"38",
          9083 => x"10",
          9084 => x"51",
          9085 => x"f4",
          9086 => x"a0",
          9087 => x"8c",
          9088 => x"58",
          9089 => x"81",
          9090 => x"77",
          9091 => x"59",
          9092 => x"55",
          9093 => x"02",
          9094 => x"33",
          9095 => x"58",
          9096 => x"2e",
          9097 => x"80",
          9098 => x"1f",
          9099 => x"94",
          9100 => x"8c",
          9101 => x"58",
          9102 => x"61",
          9103 => x"77",
          9104 => x"59",
          9105 => x"81",
          9106 => x"ff",
          9107 => x"ef",
          9108 => x"27",
          9109 => x"7a",
          9110 => x"57",
          9111 => x"b8",
          9112 => x"1a",
          9113 => x"58",
          9114 => x"77",
          9115 => x"81",
          9116 => x"ff",
          9117 => x"90",
          9118 => x"44",
          9119 => x"60",
          9120 => x"38",
          9121 => x"a1",
          9122 => x"18",
          9123 => x"25",
          9124 => x"22",
          9125 => x"38",
          9126 => x"05",
          9127 => x"57",
          9128 => x"07",
          9129 => x"b9",
          9130 => x"38",
          9131 => x"74",
          9132 => x"16",
          9133 => x"84",
          9134 => x"56",
          9135 => x"77",
          9136 => x"fe",
          9137 => x"7a",
          9138 => x"78",
          9139 => x"79",
          9140 => x"a0",
          9141 => x"81",
          9142 => x"78",
          9143 => x"38",
          9144 => x"33",
          9145 => x"a0",
          9146 => x"06",
          9147 => x"16",
          9148 => x"77",
          9149 => x"38",
          9150 => x"05",
          9151 => x"19",
          9152 => x"59",
          9153 => x"34",
          9154 => x"87",
          9155 => x"51",
          9156 => x"84",
          9157 => x"8b",
          9158 => x"5b",
          9159 => x"27",
          9160 => x"87",
          9161 => x"e4",
          9162 => x"38",
          9163 => x"08",
          9164 => x"e4",
          9165 => x"09",
          9166 => x"d6",
          9167 => x"db",
          9168 => x"1f",
          9169 => x"02",
          9170 => x"db",
          9171 => x"58",
          9172 => x"81",
          9173 => x"5b",
          9174 => x"90",
          9175 => x"8c",
          9176 => x"8a",
          9177 => x"b8",
          9178 => x"5b",
          9179 => x"51",
          9180 => x"84",
          9181 => x"56",
          9182 => x"08",
          9183 => x"84",
          9184 => x"b8",
          9185 => x"98",
          9186 => x"80",
          9187 => x"08",
          9188 => x"f3",
          9189 => x"33",
          9190 => x"2e",
          9191 => x"82",
          9192 => x"54",
          9193 => x"18",
          9194 => x"33",
          9195 => x"3f",
          9196 => x"08",
          9197 => x"38",
          9198 => x"57",
          9199 => x"0c",
          9200 => x"bc",
          9201 => x"08",
          9202 => x"42",
          9203 => x"2e",
          9204 => x"74",
          9205 => x"25",
          9206 => x"5f",
          9207 => x"81",
          9208 => x"19",
          9209 => x"2e",
          9210 => x"81",
          9211 => x"ee",
          9212 => x"b8",
          9213 => x"84",
          9214 => x"80",
          9215 => x"38",
          9216 => x"84",
          9217 => x"38",
          9218 => x"81",
          9219 => x"1b",
          9220 => x"f3",
          9221 => x"08",
          9222 => x"08",
          9223 => x"38",
          9224 => x"78",
          9225 => x"84",
          9226 => x"54",
          9227 => x"1c",
          9228 => x"33",
          9229 => x"3f",
          9230 => x"08",
          9231 => x"38",
          9232 => x"56",
          9233 => x"0c",
          9234 => x"80",
          9235 => x"0b",
          9236 => x"57",
          9237 => x"70",
          9238 => x"34",
          9239 => x"74",
          9240 => x"0b",
          9241 => x"7b",
          9242 => x"75",
          9243 => x"57",
          9244 => x"81",
          9245 => x"ff",
          9246 => x"ef",
          9247 => x"08",
          9248 => x"98",
          9249 => x"7c",
          9250 => x"81",
          9251 => x"34",
          9252 => x"84",
          9253 => x"98",
          9254 => x"81",
          9255 => x"80",
          9256 => x"57",
          9257 => x"fe",
          9258 => x"59",
          9259 => x"51",
          9260 => x"84",
          9261 => x"56",
          9262 => x"08",
          9263 => x"c7",
          9264 => x"39",
          9265 => x"18",
          9266 => x"52",
          9267 => x"51",
          9268 => x"84",
          9269 => x"77",
          9270 => x"06",
          9271 => x"84",
          9272 => x"83",
          9273 => x"18",
          9274 => x"08",
          9275 => x"a0",
          9276 => x"8b",
          9277 => x"33",
          9278 => x"2e",
          9279 => x"84",
          9280 => x"57",
          9281 => x"7f",
          9282 => x"1f",
          9283 => x"53",
          9284 => x"e9",
          9285 => x"b8",
          9286 => x"84",
          9287 => x"fe",
          9288 => x"84",
          9289 => x"56",
          9290 => x"74",
          9291 => x"81",
          9292 => x"78",
          9293 => x"5a",
          9294 => x"05",
          9295 => x"06",
          9296 => x"56",
          9297 => x"38",
          9298 => x"06",
          9299 => x"41",
          9300 => x"57",
          9301 => x"1c",
          9302 => x"b2",
          9303 => x"33",
          9304 => x"2e",
          9305 => x"82",
          9306 => x"54",
          9307 => x"1c",
          9308 => x"33",
          9309 => x"3f",
          9310 => x"08",
          9311 => x"38",
          9312 => x"56",
          9313 => x"0c",
          9314 => x"fe",
          9315 => x"1c",
          9316 => x"08",
          9317 => x"06",
          9318 => x"60",
          9319 => x"8f",
          9320 => x"34",
          9321 => x"34",
          9322 => x"34",
          9323 => x"34",
          9324 => x"f3",
          9325 => x"5a",
          9326 => x"83",
          9327 => x"8b",
          9328 => x"1f",
          9329 => x"1b",
          9330 => x"83",
          9331 => x"33",
          9332 => x"76",
          9333 => x"05",
          9334 => x"88",
          9335 => x"75",
          9336 => x"38",
          9337 => x"57",
          9338 => x"8c",
          9339 => x"38",
          9340 => x"ff",
          9341 => x"38",
          9342 => x"70",
          9343 => x"76",
          9344 => x"a6",
          9345 => x"34",
          9346 => x"1d",
          9347 => x"7d",
          9348 => x"3f",
          9349 => x"08",
          9350 => x"e4",
          9351 => x"38",
          9352 => x"40",
          9353 => x"38",
          9354 => x"81",
          9355 => x"08",
          9356 => x"70",
          9357 => x"33",
          9358 => x"96",
          9359 => x"84",
          9360 => x"fc",
          9361 => x"b8",
          9362 => x"1d",
          9363 => x"08",
          9364 => x"31",
          9365 => x"08",
          9366 => x"a0",
          9367 => x"fb",
          9368 => x"1c",
          9369 => x"82",
          9370 => x"06",
          9371 => x"81",
          9372 => x"08",
          9373 => x"05",
          9374 => x"81",
          9375 => x"cf",
          9376 => x"56",
          9377 => x"76",
          9378 => x"70",
          9379 => x"56",
          9380 => x"2e",
          9381 => x"fa",
          9382 => x"ff",
          9383 => x"57",
          9384 => x"2e",
          9385 => x"fa",
          9386 => x"80",
          9387 => x"fe",
          9388 => x"54",
          9389 => x"53",
          9390 => x"1c",
          9391 => x"92",
          9392 => x"e4",
          9393 => x"09",
          9394 => x"38",
          9395 => x"08",
          9396 => x"b4",
          9397 => x"1d",
          9398 => x"74",
          9399 => x"27",
          9400 => x"1c",
          9401 => x"82",
          9402 => x"84",
          9403 => x"56",
          9404 => x"75",
          9405 => x"58",
          9406 => x"fa",
          9407 => x"87",
          9408 => x"57",
          9409 => x"81",
          9410 => x"75",
          9411 => x"fe",
          9412 => x"39",
          9413 => x"1c",
          9414 => x"08",
          9415 => x"52",
          9416 => x"51",
          9417 => x"fc",
          9418 => x"54",
          9419 => x"a0",
          9420 => x"53",
          9421 => x"18",
          9422 => x"96",
          9423 => x"39",
          9424 => x"7f",
          9425 => x"40",
          9426 => x"0b",
          9427 => x"98",
          9428 => x"2e",
          9429 => x"ac",
          9430 => x"2e",
          9431 => x"80",
          9432 => x"8c",
          9433 => x"22",
          9434 => x"5c",
          9435 => x"2e",
          9436 => x"54",
          9437 => x"22",
          9438 => x"55",
          9439 => x"95",
          9440 => x"80",
          9441 => x"ff",
          9442 => x"5a",
          9443 => x"26",
          9444 => x"73",
          9445 => x"11",
          9446 => x"58",
          9447 => x"d4",
          9448 => x"70",
          9449 => x"30",
          9450 => x"5c",
          9451 => x"94",
          9452 => x"0b",
          9453 => x"80",
          9454 => x"59",
          9455 => x"1c",
          9456 => x"33",
          9457 => x"56",
          9458 => x"2e",
          9459 => x"85",
          9460 => x"38",
          9461 => x"70",
          9462 => x"07",
          9463 => x"5b",
          9464 => x"26",
          9465 => x"80",
          9466 => x"ae",
          9467 => x"05",
          9468 => x"18",
          9469 => x"70",
          9470 => x"34",
          9471 => x"8a",
          9472 => x"ba",
          9473 => x"88",
          9474 => x"0b",
          9475 => x"96",
          9476 => x"72",
          9477 => x"81",
          9478 => x"0b",
          9479 => x"81",
          9480 => x"94",
          9481 => x"0b",
          9482 => x"9c",
          9483 => x"11",
          9484 => x"73",
          9485 => x"89",
          9486 => x"1c",
          9487 => x"13",
          9488 => x"34",
          9489 => x"9c",
          9490 => x"33",
          9491 => x"71",
          9492 => x"88",
          9493 => x"14",
          9494 => x"07",
          9495 => x"33",
          9496 => x"0c",
          9497 => x"33",
          9498 => x"71",
          9499 => x"5f",
          9500 => x"5a",
          9501 => x"77",
          9502 => x"99",
          9503 => x"16",
          9504 => x"2b",
          9505 => x"7b",
          9506 => x"8f",
          9507 => x"81",
          9508 => x"c0",
          9509 => x"96",
          9510 => x"7a",
          9511 => x"57",
          9512 => x"7a",
          9513 => x"07",
          9514 => x"89",
          9515 => x"e4",
          9516 => x"ff",
          9517 => x"ff",
          9518 => x"38",
          9519 => x"81",
          9520 => x"88",
          9521 => x"7a",
          9522 => x"18",
          9523 => x"05",
          9524 => x"8c",
          9525 => x"5b",
          9526 => x"11",
          9527 => x"57",
          9528 => x"90",
          9529 => x"39",
          9530 => x"30",
          9531 => x"80",
          9532 => x"25",
          9533 => x"57",
          9534 => x"38",
          9535 => x"81",
          9536 => x"80",
          9537 => x"08",
          9538 => x"39",
          9539 => x"1f",
          9540 => x"57",
          9541 => x"fe",
          9542 => x"96",
          9543 => x"59",
          9544 => x"33",
          9545 => x"5a",
          9546 => x"26",
          9547 => x"1c",
          9548 => x"33",
          9549 => x"76",
          9550 => x"72",
          9551 => x"72",
          9552 => x"7d",
          9553 => x"38",
          9554 => x"83",
          9555 => x"55",
          9556 => x"70",
          9557 => x"34",
          9558 => x"16",
          9559 => x"89",
          9560 => x"57",
          9561 => x"79",
          9562 => x"fd",
          9563 => x"83",
          9564 => x"39",
          9565 => x"70",
          9566 => x"30",
          9567 => x"5d",
          9568 => x"a9",
          9569 => x"0d",
          9570 => x"70",
          9571 => x"80",
          9572 => x"57",
          9573 => x"af",
          9574 => x"81",
          9575 => x"dc",
          9576 => x"38",
          9577 => x"81",
          9578 => x"16",
          9579 => x"0c",
          9580 => x"3d",
          9581 => x"42",
          9582 => x"27",
          9583 => x"73",
          9584 => x"08",
          9585 => x"61",
          9586 => x"05",
          9587 => x"53",
          9588 => x"38",
          9589 => x"73",
          9590 => x"ec",
          9591 => x"ff",
          9592 => x"38",
          9593 => x"56",
          9594 => x"81",
          9595 => x"83",
          9596 => x"70",
          9597 => x"30",
          9598 => x"71",
          9599 => x"57",
          9600 => x"73",
          9601 => x"74",
          9602 => x"82",
          9603 => x"80",
          9604 => x"38",
          9605 => x"0b",
          9606 => x"33",
          9607 => x"06",
          9608 => x"73",
          9609 => x"ab",
          9610 => x"2e",
          9611 => x"16",
          9612 => x"81",
          9613 => x"54",
          9614 => x"38",
          9615 => x"06",
          9616 => x"84",
          9617 => x"fe",
          9618 => x"38",
          9619 => x"5d",
          9620 => x"81",
          9621 => x"70",
          9622 => x"33",
          9623 => x"73",
          9624 => x"f0",
          9625 => x"39",
          9626 => x"dc",
          9627 => x"70",
          9628 => x"07",
          9629 => x"55",
          9630 => x"a1",
          9631 => x"70",
          9632 => x"74",
          9633 => x"72",
          9634 => x"38",
          9635 => x"32",
          9636 => x"80",
          9637 => x"51",
          9638 => x"e1",
          9639 => x"1d",
          9640 => x"96",
          9641 => x"41",
          9642 => x"9f",
          9643 => x"38",
          9644 => x"b5",
          9645 => x"81",
          9646 => x"84",
          9647 => x"83",
          9648 => x"54",
          9649 => x"38",
          9650 => x"84",
          9651 => x"93",
          9652 => x"83",
          9653 => x"70",
          9654 => x"5c",
          9655 => x"2e",
          9656 => x"e4",
          9657 => x"0b",
          9658 => x"80",
          9659 => x"de",
          9660 => x"b8",
          9661 => x"b8",
          9662 => x"3d",
          9663 => x"73",
          9664 => x"70",
          9665 => x"25",
          9666 => x"55",
          9667 => x"80",
          9668 => x"81",
          9669 => x"62",
          9670 => x"55",
          9671 => x"2e",
          9672 => x"80",
          9673 => x"30",
          9674 => x"78",
          9675 => x"59",
          9676 => x"73",
          9677 => x"75",
          9678 => x"5a",
          9679 => x"84",
          9680 => x"82",
          9681 => x"38",
          9682 => x"76",
          9683 => x"38",
          9684 => x"11",
          9685 => x"22",
          9686 => x"70",
          9687 => x"2a",
          9688 => x"5f",
          9689 => x"ae",
          9690 => x"72",
          9691 => x"17",
          9692 => x"38",
          9693 => x"19",
          9694 => x"23",
          9695 => x"fe",
          9696 => x"78",
          9697 => x"ff",
          9698 => x"58",
          9699 => x"7a",
          9700 => x"e6",
          9701 => x"ff",
          9702 => x"72",
          9703 => x"f1",
          9704 => x"2e",
          9705 => x"19",
          9706 => x"22",
          9707 => x"ae",
          9708 => x"76",
          9709 => x"05",
          9710 => x"57",
          9711 => x"8f",
          9712 => x"70",
          9713 => x"7c",
          9714 => x"81",
          9715 => x"8b",
          9716 => x"55",
          9717 => x"70",
          9718 => x"34",
          9719 => x"72",
          9720 => x"73",
          9721 => x"78",
          9722 => x"81",
          9723 => x"54",
          9724 => x"2e",
          9725 => x"74",
          9726 => x"d0",
          9727 => x"32",
          9728 => x"80",
          9729 => x"54",
          9730 => x"85",
          9731 => x"83",
          9732 => x"59",
          9733 => x"83",
          9734 => x"75",
          9735 => x"30",
          9736 => x"80",
          9737 => x"07",
          9738 => x"54",
          9739 => x"83",
          9740 => x"8b",
          9741 => x"38",
          9742 => x"8a",
          9743 => x"07",
          9744 => x"26",
          9745 => x"56",
          9746 => x"7e",
          9747 => x"fc",
          9748 => x"57",
          9749 => x"15",
          9750 => x"18",
          9751 => x"74",
          9752 => x"a0",
          9753 => x"76",
          9754 => x"83",
          9755 => x"88",
          9756 => x"38",
          9757 => x"58",
          9758 => x"82",
          9759 => x"83",
          9760 => x"83",
          9761 => x"38",
          9762 => x"81",
          9763 => x"9d",
          9764 => x"06",
          9765 => x"2e",
          9766 => x"90",
          9767 => x"82",
          9768 => x"5e",
          9769 => x"85",
          9770 => x"07",
          9771 => x"1d",
          9772 => x"e4",
          9773 => x"b8",
          9774 => x"1d",
          9775 => x"84",
          9776 => x"80",
          9777 => x"38",
          9778 => x"08",
          9779 => x"81",
          9780 => x"38",
          9781 => x"81",
          9782 => x"80",
          9783 => x"38",
          9784 => x"81",
          9785 => x"82",
          9786 => x"08",
          9787 => x"73",
          9788 => x"08",
          9789 => x"f9",
          9790 => x"16",
          9791 => x"11",
          9792 => x"40",
          9793 => x"a0",
          9794 => x"75",
          9795 => x"85",
          9796 => x"07",
          9797 => x"39",
          9798 => x"56",
          9799 => x"09",
          9800 => x"ac",
          9801 => x"54",
          9802 => x"09",
          9803 => x"a0",
          9804 => x"18",
          9805 => x"23",
          9806 => x"1d",
          9807 => x"54",
          9808 => x"83",
          9809 => x"73",
          9810 => x"05",
          9811 => x"13",
          9812 => x"27",
          9813 => x"a0",
          9814 => x"ab",
          9815 => x"51",
          9816 => x"84",
          9817 => x"ab",
          9818 => x"54",
          9819 => x"08",
          9820 => x"74",
          9821 => x"06",
          9822 => x"ce",
          9823 => x"33",
          9824 => x"81",
          9825 => x"74",
          9826 => x"cd",
          9827 => x"08",
          9828 => x"60",
          9829 => x"11",
          9830 => x"12",
          9831 => x"2b",
          9832 => x"41",
          9833 => x"7d",
          9834 => x"d8",
          9835 => x"1d",
          9836 => x"65",
          9837 => x"b7",
          9838 => x"55",
          9839 => x"fe",
          9840 => x"17",
          9841 => x"88",
          9842 => x"39",
          9843 => x"76",
          9844 => x"fd",
          9845 => x"82",
          9846 => x"06",
          9847 => x"59",
          9848 => x"2e",
          9849 => x"fd",
          9850 => x"82",
          9851 => x"98",
          9852 => x"a0",
          9853 => x"88",
          9854 => x"06",
          9855 => x"d6",
          9856 => x"0b",
          9857 => x"80",
          9858 => x"e4",
          9859 => x"0d",
          9860 => x"ff",
          9861 => x"81",
          9862 => x"80",
          9863 => x"1d",
          9864 => x"26",
          9865 => x"79",
          9866 => x"77",
          9867 => x"5a",
          9868 => x"79",
          9869 => x"83",
          9870 => x"51",
          9871 => x"3f",
          9872 => x"08",
          9873 => x"06",
          9874 => x"81",
          9875 => x"78",
          9876 => x"38",
          9877 => x"06",
          9878 => x"11",
          9879 => x"74",
          9880 => x"ff",
          9881 => x"80",
          9882 => x"38",
          9883 => x"0b",
          9884 => x"33",
          9885 => x"06",
          9886 => x"73",
          9887 => x"e0",
          9888 => x"2e",
          9889 => x"19",
          9890 => x"81",
          9891 => x"54",
          9892 => x"38",
          9893 => x"06",
          9894 => x"d4",
          9895 => x"15",
          9896 => x"26",
          9897 => x"82",
          9898 => x"ff",
          9899 => x"ff",
          9900 => x"78",
          9901 => x"38",
          9902 => x"70",
          9903 => x"e0",
          9904 => x"ff",
          9905 => x"56",
          9906 => x"1b",
          9907 => x"74",
          9908 => x"1b",
          9909 => x"55",
          9910 => x"80",
          9911 => x"39",
          9912 => x"33",
          9913 => x"06",
          9914 => x"80",
          9915 => x"38",
          9916 => x"83",
          9917 => x"a0",
          9918 => x"55",
          9919 => x"81",
          9920 => x"39",
          9921 => x"33",
          9922 => x"33",
          9923 => x"71",
          9924 => x"77",
          9925 => x"0c",
          9926 => x"95",
          9927 => x"a0",
          9928 => x"2a",
          9929 => x"74",
          9930 => x"7c",
          9931 => x"5a",
          9932 => x"34",
          9933 => x"ff",
          9934 => x"83",
          9935 => x"33",
          9936 => x"81",
          9937 => x"81",
          9938 => x"38",
          9939 => x"74",
          9940 => x"06",
          9941 => x"f2",
          9942 => x"84",
          9943 => x"93",
          9944 => x"eb",
          9945 => x"69",
          9946 => x"80",
          9947 => x"42",
          9948 => x"61",
          9949 => x"08",
          9950 => x"42",
          9951 => x"85",
          9952 => x"70",
          9953 => x"33",
          9954 => x"56",
          9955 => x"2e",
          9956 => x"74",
          9957 => x"ba",
          9958 => x"38",
          9959 => x"33",
          9960 => x"24",
          9961 => x"75",
          9962 => x"d0",
          9963 => x"08",
          9964 => x"58",
          9965 => x"85",
          9966 => x"61",
          9967 => x"fe",
          9968 => x"5d",
          9969 => x"2e",
          9970 => x"17",
          9971 => x"bb",
          9972 => x"b8",
          9973 => x"ff",
          9974 => x"06",
          9975 => x"80",
          9976 => x"38",
          9977 => x"75",
          9978 => x"b8",
          9979 => x"81",
          9980 => x"52",
          9981 => x"51",
          9982 => x"3f",
          9983 => x"08",
          9984 => x"70",
          9985 => x"56",
          9986 => x"84",
          9987 => x"80",
          9988 => x"75",
          9989 => x"06",
          9990 => x"60",
          9991 => x"80",
          9992 => x"18",
          9993 => x"b4",
          9994 => x"7b",
          9995 => x"54",
          9996 => x"17",
          9997 => x"18",
          9998 => x"ff",
          9999 => x"84",
         10000 => x"7b",
         10001 => x"ff",
         10002 => x"74",
         10003 => x"84",
         10004 => x"38",
         10005 => x"33",
         10006 => x"33",
         10007 => x"07",
         10008 => x"56",
         10009 => x"d5",
         10010 => x"38",
         10011 => x"8b",
         10012 => x"d9",
         10013 => x"61",
         10014 => x"81",
         10015 => x"2e",
         10016 => x"8d",
         10017 => x"26",
         10018 => x"80",
         10019 => x"80",
         10020 => x"71",
         10021 => x"5e",
         10022 => x"80",
         10023 => x"06",
         10024 => x"80",
         10025 => x"80",
         10026 => x"71",
         10027 => x"57",
         10028 => x"38",
         10029 => x"83",
         10030 => x"12",
         10031 => x"2b",
         10032 => x"07",
         10033 => x"70",
         10034 => x"2b",
         10035 => x"07",
         10036 => x"43",
         10037 => x"75",
         10038 => x"80",
         10039 => x"82",
         10040 => x"c8",
         10041 => x"11",
         10042 => x"06",
         10043 => x"8d",
         10044 => x"26",
         10045 => x"78",
         10046 => x"76",
         10047 => x"c5",
         10048 => x"5f",
         10049 => x"18",
         10050 => x"77",
         10051 => x"c4",
         10052 => x"78",
         10053 => x"87",
         10054 => x"ca",
         10055 => x"c9",
         10056 => x"88",
         10057 => x"40",
         10058 => x"23",
         10059 => x"06",
         10060 => x"58",
         10061 => x"38",
         10062 => x"33",
         10063 => x"33",
         10064 => x"07",
         10065 => x"a4",
         10066 => x"17",
         10067 => x"82",
         10068 => x"90",
         10069 => x"2b",
         10070 => x"33",
         10071 => x"88",
         10072 => x"71",
         10073 => x"5a",
         10074 => x"42",
         10075 => x"33",
         10076 => x"33",
         10077 => x"07",
         10078 => x"58",
         10079 => x"81",
         10080 => x"1c",
         10081 => x"05",
         10082 => x"26",
         10083 => x"78",
         10084 => x"31",
         10085 => x"8e",
         10086 => x"e4",
         10087 => x"b8",
         10088 => x"2e",
         10089 => x"84",
         10090 => x"80",
         10091 => x"f5",
         10092 => x"83",
         10093 => x"ff",
         10094 => x"38",
         10095 => x"9f",
         10096 => x"eb",
         10097 => x"82",
         10098 => x"19",
         10099 => x"19",
         10100 => x"70",
         10101 => x"7b",
         10102 => x"0c",
         10103 => x"83",
         10104 => x"38",
         10105 => x"5c",
         10106 => x"80",
         10107 => x"38",
         10108 => x"18",
         10109 => x"55",
         10110 => x"8d",
         10111 => x"19",
         10112 => x"7a",
         10113 => x"56",
         10114 => x"15",
         10115 => x"8d",
         10116 => x"18",
         10117 => x"38",
         10118 => x"18",
         10119 => x"90",
         10120 => x"80",
         10121 => x"34",
         10122 => x"86",
         10123 => x"77",
         10124 => x"bc",
         10125 => x"5d",
         10126 => x"bc",
         10127 => x"18",
         10128 => x"c4",
         10129 => x"0c",
         10130 => x"18",
         10131 => x"77",
         10132 => x"0c",
         10133 => x"04",
         10134 => x"b8",
         10135 => x"3d",
         10136 => x"33",
         10137 => x"81",
         10138 => x"57",
         10139 => x"26",
         10140 => x"17",
         10141 => x"06",
         10142 => x"59",
         10143 => x"87",
         10144 => x"7e",
         10145 => x"d4",
         10146 => x"7c",
         10147 => x"5b",
         10148 => x"05",
         10149 => x"70",
         10150 => x"33",
         10151 => x"5a",
         10152 => x"99",
         10153 => x"e0",
         10154 => x"ff",
         10155 => x"ff",
         10156 => x"77",
         10157 => x"38",
         10158 => x"81",
         10159 => x"55",
         10160 => x"9f",
         10161 => x"75",
         10162 => x"81",
         10163 => x"77",
         10164 => x"78",
         10165 => x"30",
         10166 => x"9f",
         10167 => x"5d",
         10168 => x"80",
         10169 => x"38",
         10170 => x"1e",
         10171 => x"7c",
         10172 => x"38",
         10173 => x"a9",
         10174 => x"2e",
         10175 => x"77",
         10176 => x"06",
         10177 => x"7d",
         10178 => x"80",
         10179 => x"39",
         10180 => x"57",
         10181 => x"e9",
         10182 => x"06",
         10183 => x"59",
         10184 => x"32",
         10185 => x"80",
         10186 => x"5a",
         10187 => x"83",
         10188 => x"81",
         10189 => x"a6",
         10190 => x"77",
         10191 => x"59",
         10192 => x"33",
         10193 => x"7a",
         10194 => x"38",
         10195 => x"33",
         10196 => x"33",
         10197 => x"71",
         10198 => x"83",
         10199 => x"70",
         10200 => x"2b",
         10201 => x"33",
         10202 => x"59",
         10203 => x"40",
         10204 => x"84",
         10205 => x"ff",
         10206 => x"57",
         10207 => x"25",
         10208 => x"84",
         10209 => x"33",
         10210 => x"9f",
         10211 => x"31",
         10212 => x"10",
         10213 => x"05",
         10214 => x"44",
         10215 => x"5b",
         10216 => x"5b",
         10217 => x"80",
         10218 => x"38",
         10219 => x"18",
         10220 => x"b4",
         10221 => x"55",
         10222 => x"ff",
         10223 => x"81",
         10224 => x"b8",
         10225 => x"17",
         10226 => x"b4",
         10227 => x"b8",
         10228 => x"2e",
         10229 => x"55",
         10230 => x"b4",
         10231 => x"58",
         10232 => x"81",
         10233 => x"33",
         10234 => x"07",
         10235 => x"58",
         10236 => x"d5",
         10237 => x"06",
         10238 => x"0b",
         10239 => x"57",
         10240 => x"e9",
         10241 => x"38",
         10242 => x"32",
         10243 => x"80",
         10244 => x"42",
         10245 => x"bc",
         10246 => x"e8",
         10247 => x"82",
         10248 => x"ff",
         10249 => x"0b",
         10250 => x"1e",
         10251 => x"7b",
         10252 => x"81",
         10253 => x"81",
         10254 => x"27",
         10255 => x"77",
         10256 => x"b7",
         10257 => x"84",
         10258 => x"83",
         10259 => x"d1",
         10260 => x"39",
         10261 => x"ee",
         10262 => x"94",
         10263 => x"7b",
         10264 => x"5d",
         10265 => x"81",
         10266 => x"71",
         10267 => x"1b",
         10268 => x"56",
         10269 => x"80",
         10270 => x"80",
         10271 => x"85",
         10272 => x"18",
         10273 => x"40",
         10274 => x"70",
         10275 => x"33",
         10276 => x"05",
         10277 => x"71",
         10278 => x"5b",
         10279 => x"77",
         10280 => x"8e",
         10281 => x"2e",
         10282 => x"58",
         10283 => x"8d",
         10284 => x"93",
         10285 => x"b8",
         10286 => x"3d",
         10287 => x"58",
         10288 => x"fe",
         10289 => x"0b",
         10290 => x"83",
         10291 => x"5d",
         10292 => x"39",
         10293 => x"b8",
         10294 => x"3d",
         10295 => x"0b",
         10296 => x"83",
         10297 => x"5a",
         10298 => x"81",
         10299 => x"7a",
         10300 => x"5c",
         10301 => x"31",
         10302 => x"57",
         10303 => x"80",
         10304 => x"38",
         10305 => x"e1",
         10306 => x"81",
         10307 => x"e4",
         10308 => x"58",
         10309 => x"05",
         10310 => x"70",
         10311 => x"33",
         10312 => x"ff",
         10313 => x"42",
         10314 => x"2e",
         10315 => x"75",
         10316 => x"38",
         10317 => x"57",
         10318 => x"fc",
         10319 => x"58",
         10320 => x"80",
         10321 => x"80",
         10322 => x"71",
         10323 => x"57",
         10324 => x"2e",
         10325 => x"f9",
         10326 => x"1b",
         10327 => x"b4",
         10328 => x"2e",
         10329 => x"17",
         10330 => x"7a",
         10331 => x"06",
         10332 => x"81",
         10333 => x"b8",
         10334 => x"17",
         10335 => x"b0",
         10336 => x"b8",
         10337 => x"2e",
         10338 => x"58",
         10339 => x"b4",
         10340 => x"f9",
         10341 => x"84",
         10342 => x"b7",
         10343 => x"b6",
         10344 => x"88",
         10345 => x"5e",
         10346 => x"d5",
         10347 => x"06",
         10348 => x"b8",
         10349 => x"33",
         10350 => x"71",
         10351 => x"88",
         10352 => x"14",
         10353 => x"07",
         10354 => x"33",
         10355 => x"41",
         10356 => x"5c",
         10357 => x"8b",
         10358 => x"2e",
         10359 => x"f8",
         10360 => x"9c",
         10361 => x"33",
         10362 => x"71",
         10363 => x"88",
         10364 => x"14",
         10365 => x"07",
         10366 => x"33",
         10367 => x"44",
         10368 => x"5a",
         10369 => x"8a",
         10370 => x"2e",
         10371 => x"f8",
         10372 => x"a0",
         10373 => x"33",
         10374 => x"71",
         10375 => x"88",
         10376 => x"14",
         10377 => x"07",
         10378 => x"33",
         10379 => x"1e",
         10380 => x"a4",
         10381 => x"33",
         10382 => x"71",
         10383 => x"88",
         10384 => x"14",
         10385 => x"07",
         10386 => x"33",
         10387 => x"90",
         10388 => x"44",
         10389 => x"45",
         10390 => x"56",
         10391 => x"34",
         10392 => x"22",
         10393 => x"7c",
         10394 => x"23",
         10395 => x"23",
         10396 => x"0b",
         10397 => x"80",
         10398 => x"0c",
         10399 => x"7b",
         10400 => x"f0",
         10401 => x"7f",
         10402 => x"95",
         10403 => x"b4",
         10404 => x"b8",
         10405 => x"81",
         10406 => x"59",
         10407 => x"3f",
         10408 => x"08",
         10409 => x"81",
         10410 => x"38",
         10411 => x"08",
         10412 => x"b4",
         10413 => x"18",
         10414 => x"7f",
         10415 => x"27",
         10416 => x"17",
         10417 => x"82",
         10418 => x"38",
         10419 => x"08",
         10420 => x"39",
         10421 => x"80",
         10422 => x"38",
         10423 => x"8a",
         10424 => x"98",
         10425 => x"fc",
         10426 => x"e3",
         10427 => x"e2",
         10428 => x"88",
         10429 => x"5a",
         10430 => x"f6",
         10431 => x"17",
         10432 => x"f6",
         10433 => x"e4",
         10434 => x"33",
         10435 => x"71",
         10436 => x"88",
         10437 => x"14",
         10438 => x"07",
         10439 => x"33",
         10440 => x"1e",
         10441 => x"82",
         10442 => x"44",
         10443 => x"f5",
         10444 => x"58",
         10445 => x"f9",
         10446 => x"58",
         10447 => x"75",
         10448 => x"a8",
         10449 => x"77",
         10450 => x"59",
         10451 => x"75",
         10452 => x"da",
         10453 => x"39",
         10454 => x"17",
         10455 => x"08",
         10456 => x"52",
         10457 => x"51",
         10458 => x"3f",
         10459 => x"f0",
         10460 => x"80",
         10461 => x"64",
         10462 => x"3d",
         10463 => x"ff",
         10464 => x"75",
         10465 => x"e9",
         10466 => x"81",
         10467 => x"70",
         10468 => x"55",
         10469 => x"80",
         10470 => x"ed",
         10471 => x"2e",
         10472 => x"84",
         10473 => x"54",
         10474 => x"80",
         10475 => x"10",
         10476 => x"ac",
         10477 => x"55",
         10478 => x"2e",
         10479 => x"74",
         10480 => x"73",
         10481 => x"38",
         10482 => x"62",
         10483 => x"0c",
         10484 => x"80",
         10485 => x"80",
         10486 => x"70",
         10487 => x"51",
         10488 => x"84",
         10489 => x"54",
         10490 => x"e4",
         10491 => x"0d",
         10492 => x"84",
         10493 => x"92",
         10494 => x"75",
         10495 => x"70",
         10496 => x"56",
         10497 => x"89",
         10498 => x"82",
         10499 => x"ff",
         10500 => x"5c",
         10501 => x"2e",
         10502 => x"80",
         10503 => x"e4",
         10504 => x"5b",
         10505 => x"59",
         10506 => x"81",
         10507 => x"78",
         10508 => x"5a",
         10509 => x"12",
         10510 => x"76",
         10511 => x"38",
         10512 => x"81",
         10513 => x"54",
         10514 => x"57",
         10515 => x"89",
         10516 => x"70",
         10517 => x"57",
         10518 => x"70",
         10519 => x"54",
         10520 => x"09",
         10521 => x"38",
         10522 => x"38",
         10523 => x"70",
         10524 => x"07",
         10525 => x"07",
         10526 => x"79",
         10527 => x"38",
         10528 => x"1d",
         10529 => x"7b",
         10530 => x"38",
         10531 => x"98",
         10532 => x"24",
         10533 => x"79",
         10534 => x"fe",
         10535 => x"3d",
         10536 => x"84",
         10537 => x"05",
         10538 => x"89",
         10539 => x"2e",
         10540 => x"bf",
         10541 => x"9d",
         10542 => x"53",
         10543 => x"05",
         10544 => x"9f",
         10545 => x"e4",
         10546 => x"b8",
         10547 => x"2e",
         10548 => x"79",
         10549 => x"75",
         10550 => x"0c",
         10551 => x"04",
         10552 => x"52",
         10553 => x"52",
         10554 => x"3f",
         10555 => x"08",
         10556 => x"e4",
         10557 => x"81",
         10558 => x"9c",
         10559 => x"80",
         10560 => x"38",
         10561 => x"83",
         10562 => x"84",
         10563 => x"38",
         10564 => x"58",
         10565 => x"38",
         10566 => x"81",
         10567 => x"80",
         10568 => x"38",
         10569 => x"33",
         10570 => x"71",
         10571 => x"61",
         10572 => x"58",
         10573 => x"7d",
         10574 => x"e9",
         10575 => x"8e",
         10576 => x"0b",
         10577 => x"a1",
         10578 => x"34",
         10579 => x"91",
         10580 => x"56",
         10581 => x"17",
         10582 => x"57",
         10583 => x"9a",
         10584 => x"0b",
         10585 => x"7d",
         10586 => x"83",
         10587 => x"38",
         10588 => x"0b",
         10589 => x"80",
         10590 => x"34",
         10591 => x"1c",
         10592 => x"9f",
         10593 => x"55",
         10594 => x"16",
         10595 => x"2e",
         10596 => x"7e",
         10597 => x"7d",
         10598 => x"57",
         10599 => x"7c",
         10600 => x"9c",
         10601 => x"26",
         10602 => x"82",
         10603 => x"0c",
         10604 => x"02",
         10605 => x"33",
         10606 => x"5d",
         10607 => x"25",
         10608 => x"86",
         10609 => x"5e",
         10610 => x"b8",
         10611 => x"82",
         10612 => x"c2",
         10613 => x"84",
         10614 => x"5d",
         10615 => x"91",
         10616 => x"2a",
         10617 => x"7d",
         10618 => x"38",
         10619 => x"5a",
         10620 => x"38",
         10621 => x"81",
         10622 => x"80",
         10623 => x"77",
         10624 => x"58",
         10625 => x"08",
         10626 => x"67",
         10627 => x"67",
         10628 => x"9a",
         10629 => x"88",
         10630 => x"33",
         10631 => x"57",
         10632 => x"2e",
         10633 => x"7a",
         10634 => x"9c",
         10635 => x"33",
         10636 => x"71",
         10637 => x"88",
         10638 => x"14",
         10639 => x"07",
         10640 => x"33",
         10641 => x"60",
         10642 => x"60",
         10643 => x"52",
         10644 => x"5d",
         10645 => x"22",
         10646 => x"77",
         10647 => x"80",
         10648 => x"34",
         10649 => x"1a",
         10650 => x"2a",
         10651 => x"74",
         10652 => x"ac",
         10653 => x"2e",
         10654 => x"75",
         10655 => x"8a",
         10656 => x"89",
         10657 => x"5b",
         10658 => x"70",
         10659 => x"25",
         10660 => x"76",
         10661 => x"38",
         10662 => x"06",
         10663 => x"80",
         10664 => x"38",
         10665 => x"51",
         10666 => x"3f",
         10667 => x"08",
         10668 => x"e4",
         10669 => x"83",
         10670 => x"84",
         10671 => x"ff",
         10672 => x"38",
         10673 => x"56",
         10674 => x"80",
         10675 => x"91",
         10676 => x"95",
         10677 => x"2a",
         10678 => x"74",
         10679 => x"b8",
         10680 => x"80",
         10681 => x"ed",
         10682 => x"80",
         10683 => x"e5",
         10684 => x"80",
         10685 => x"dd",
         10686 => x"cd",
         10687 => x"b8",
         10688 => x"88",
         10689 => x"76",
         10690 => x"fc",
         10691 => x"76",
         10692 => x"57",
         10693 => x"95",
         10694 => x"17",
         10695 => x"2b",
         10696 => x"07",
         10697 => x"5e",
         10698 => x"39",
         10699 => x"7b",
         10700 => x"38",
         10701 => x"51",
         10702 => x"3f",
         10703 => x"08",
         10704 => x"e4",
         10705 => x"81",
         10706 => x"b8",
         10707 => x"2e",
         10708 => x"84",
         10709 => x"ff",
         10710 => x"38",
         10711 => x"52",
         10712 => x"b2",
         10713 => x"b8",
         10714 => x"90",
         10715 => x"08",
         10716 => x"19",
         10717 => x"5b",
         10718 => x"ff",
         10719 => x"16",
         10720 => x"84",
         10721 => x"07",
         10722 => x"18",
         10723 => x"7a",
         10724 => x"a0",
         10725 => x"39",
         10726 => x"17",
         10727 => x"95",
         10728 => x"cc",
         10729 => x"33",
         10730 => x"71",
         10731 => x"90",
         10732 => x"07",
         10733 => x"80",
         10734 => x"34",
         10735 => x"17",
         10736 => x"90",
         10737 => x"cc",
         10738 => x"34",
         10739 => x"0b",
         10740 => x"7e",
         10741 => x"80",
         10742 => x"34",
         10743 => x"17",
         10744 => x"5d",
         10745 => x"09",
         10746 => x"84",
         10747 => x"39",
         10748 => x"72",
         10749 => x"5d",
         10750 => x"7e",
         10751 => x"83",
         10752 => x"79",
         10753 => x"81",
         10754 => x"81",
         10755 => x"b8",
         10756 => x"16",
         10757 => x"a3",
         10758 => x"b8",
         10759 => x"2e",
         10760 => x"57",
         10761 => x"b4",
         10762 => x"56",
         10763 => x"90",
         10764 => x"7a",
         10765 => x"bc",
         10766 => x"0c",
         10767 => x"81",
         10768 => x"08",
         10769 => x"70",
         10770 => x"33",
         10771 => x"a4",
         10772 => x"b8",
         10773 => x"2e",
         10774 => x"81",
         10775 => x"b8",
         10776 => x"17",
         10777 => x"08",
         10778 => x"31",
         10779 => x"08",
         10780 => x"a0",
         10781 => x"ff",
         10782 => x"16",
         10783 => x"82",
         10784 => x"06",
         10785 => x"81",
         10786 => x"08",
         10787 => x"05",
         10788 => x"81",
         10789 => x"ff",
         10790 => x"7c",
         10791 => x"39",
         10792 => x"0c",
         10793 => x"af",
         10794 => x"1a",
         10795 => x"a2",
         10796 => x"ff",
         10797 => x"80",
         10798 => x"38",
         10799 => x"9c",
         10800 => x"05",
         10801 => x"77",
         10802 => x"df",
         10803 => x"22",
         10804 => x"b0",
         10805 => x"56",
         10806 => x"2e",
         10807 => x"75",
         10808 => x"9c",
         10809 => x"56",
         10810 => x"75",
         10811 => x"76",
         10812 => x"39",
         10813 => x"79",
         10814 => x"39",
         10815 => x"08",
         10816 => x"0c",
         10817 => x"81",
         10818 => x"fe",
         10819 => x"3d",
         10820 => x"67",
         10821 => x"5d",
         10822 => x"0c",
         10823 => x"80",
         10824 => x"79",
         10825 => x"80",
         10826 => x"75",
         10827 => x"80",
         10828 => x"86",
         10829 => x"1b",
         10830 => x"78",
         10831 => x"b7",
         10832 => x"74",
         10833 => x"76",
         10834 => x"91",
         10835 => x"74",
         10836 => x"90",
         10837 => x"06",
         10838 => x"76",
         10839 => x"ed",
         10840 => x"08",
         10841 => x"71",
         10842 => x"7b",
         10843 => x"ef",
         10844 => x"2e",
         10845 => x"60",
         10846 => x"ff",
         10847 => x"81",
         10848 => x"19",
         10849 => x"76",
         10850 => x"5b",
         10851 => x"75",
         10852 => x"88",
         10853 => x"81",
         10854 => x"85",
         10855 => x"2e",
         10856 => x"74",
         10857 => x"60",
         10858 => x"08",
         10859 => x"1a",
         10860 => x"41",
         10861 => x"27",
         10862 => x"8a",
         10863 => x"78",
         10864 => x"08",
         10865 => x"74",
         10866 => x"d5",
         10867 => x"7c",
         10868 => x"57",
         10869 => x"83",
         10870 => x"1b",
         10871 => x"27",
         10872 => x"7b",
         10873 => x"54",
         10874 => x"52",
         10875 => x"51",
         10876 => x"3f",
         10877 => x"08",
         10878 => x"60",
         10879 => x"57",
         10880 => x"2e",
         10881 => x"19",
         10882 => x"56",
         10883 => x"9e",
         10884 => x"76",
         10885 => x"b8",
         10886 => x"55",
         10887 => x"05",
         10888 => x"70",
         10889 => x"34",
         10890 => x"74",
         10891 => x"89",
         10892 => x"78",
         10893 => x"19",
         10894 => x"1e",
         10895 => x"1a",
         10896 => x"1d",
         10897 => x"7b",
         10898 => x"80",
         10899 => x"b8",
         10900 => x"3d",
         10901 => x"84",
         10902 => x"92",
         10903 => x"74",
         10904 => x"39",
         10905 => x"57",
         10906 => x"06",
         10907 => x"31",
         10908 => x"78",
         10909 => x"7b",
         10910 => x"b4",
         10911 => x"2e",
         10912 => x"0b",
         10913 => x"71",
         10914 => x"7f",
         10915 => x"81",
         10916 => x"38",
         10917 => x"53",
         10918 => x"81",
         10919 => x"ff",
         10920 => x"84",
         10921 => x"80",
         10922 => x"ff",
         10923 => x"75",
         10924 => x"7a",
         10925 => x"60",
         10926 => x"83",
         10927 => x"79",
         10928 => x"b8",
         10929 => x"77",
         10930 => x"e6",
         10931 => x"81",
         10932 => x"77",
         10933 => x"59",
         10934 => x"56",
         10935 => x"fe",
         10936 => x"70",
         10937 => x"33",
         10938 => x"05",
         10939 => x"16",
         10940 => x"38",
         10941 => x"81",
         10942 => x"08",
         10943 => x"70",
         10944 => x"33",
         10945 => x"9e",
         10946 => x"5b",
         10947 => x"08",
         10948 => x"81",
         10949 => x"38",
         10950 => x"08",
         10951 => x"b4",
         10952 => x"1a",
         10953 => x"b8",
         10954 => x"55",
         10955 => x"08",
         10956 => x"38",
         10957 => x"55",
         10958 => x"09",
         10959 => x"d4",
         10960 => x"b4",
         10961 => x"1a",
         10962 => x"7f",
         10963 => x"33",
         10964 => x"fe",
         10965 => x"fe",
         10966 => x"9c",
         10967 => x"1a",
         10968 => x"84",
         10969 => x"08",
         10970 => x"ff",
         10971 => x"84",
         10972 => x"55",
         10973 => x"81",
         10974 => x"ff",
         10975 => x"84",
         10976 => x"81",
         10977 => x"fb",
         10978 => x"7a",
         10979 => x"fb",
         10980 => x"0b",
         10981 => x"81",
         10982 => x"e4",
         10983 => x"0d",
         10984 => x"91",
         10985 => x"0b",
         10986 => x"0c",
         10987 => x"04",
         10988 => x"62",
         10989 => x"40",
         10990 => x"80",
         10991 => x"57",
         10992 => x"9f",
         10993 => x"56",
         10994 => x"97",
         10995 => x"55",
         10996 => x"8f",
         10997 => x"22",
         10998 => x"59",
         10999 => x"2e",
         11000 => x"80",
         11001 => x"76",
         11002 => x"c4",
         11003 => x"33",
         11004 => x"bc",
         11005 => x"33",
         11006 => x"81",
         11007 => x"87",
         11008 => x"2e",
         11009 => x"94",
         11010 => x"11",
         11011 => x"77",
         11012 => x"76",
         11013 => x"80",
         11014 => x"38",
         11015 => x"06",
         11016 => x"a2",
         11017 => x"11",
         11018 => x"78",
         11019 => x"5a",
         11020 => x"38",
         11021 => x"38",
         11022 => x"55",
         11023 => x"84",
         11024 => x"81",
         11025 => x"38",
         11026 => x"86",
         11027 => x"98",
         11028 => x"1a",
         11029 => x"74",
         11030 => x"60",
         11031 => x"08",
         11032 => x"2e",
         11033 => x"98",
         11034 => x"05",
         11035 => x"fe",
         11036 => x"77",
         11037 => x"f0",
         11038 => x"22",
         11039 => x"b0",
         11040 => x"56",
         11041 => x"2e",
         11042 => x"78",
         11043 => x"2a",
         11044 => x"80",
         11045 => x"38",
         11046 => x"76",
         11047 => x"38",
         11048 => x"58",
         11049 => x"53",
         11050 => x"16",
         11051 => x"9b",
         11052 => x"b8",
         11053 => x"a1",
         11054 => x"11",
         11055 => x"56",
         11056 => x"27",
         11057 => x"80",
         11058 => x"76",
         11059 => x"57",
         11060 => x"70",
         11061 => x"33",
         11062 => x"05",
         11063 => x"16",
         11064 => x"38",
         11065 => x"83",
         11066 => x"89",
         11067 => x"79",
         11068 => x"1a",
         11069 => x"1e",
         11070 => x"1b",
         11071 => x"1f",
         11072 => x"08",
         11073 => x"5e",
         11074 => x"27",
         11075 => x"56",
         11076 => x"0c",
         11077 => x"38",
         11078 => x"58",
         11079 => x"07",
         11080 => x"1b",
         11081 => x"75",
         11082 => x"0c",
         11083 => x"04",
         11084 => x"e4",
         11085 => x"0d",
         11086 => x"33",
         11087 => x"c8",
         11088 => x"fe",
         11089 => x"9c",
         11090 => x"56",
         11091 => x"06",
         11092 => x"31",
         11093 => x"79",
         11094 => x"7a",
         11095 => x"b4",
         11096 => x"2e",
         11097 => x"0b",
         11098 => x"71",
         11099 => x"7f",
         11100 => x"81",
         11101 => x"38",
         11102 => x"53",
         11103 => x"81",
         11104 => x"ff",
         11105 => x"84",
         11106 => x"80",
         11107 => x"ff",
         11108 => x"76",
         11109 => x"7b",
         11110 => x"60",
         11111 => x"83",
         11112 => x"7a",
         11113 => x"7e",
         11114 => x"78",
         11115 => x"38",
         11116 => x"05",
         11117 => x"70",
         11118 => x"34",
         11119 => x"75",
         11120 => x"58",
         11121 => x"19",
         11122 => x"39",
         11123 => x"16",
         11124 => x"16",
         11125 => x"17",
         11126 => x"ff",
         11127 => x"81",
         11128 => x"e4",
         11129 => x"09",
         11130 => x"ab",
         11131 => x"e4",
         11132 => x"34",
         11133 => x"a8",
         11134 => x"84",
         11135 => x"5d",
         11136 => x"17",
         11137 => x"f0",
         11138 => x"33",
         11139 => x"2e",
         11140 => x"fe",
         11141 => x"54",
         11142 => x"a0",
         11143 => x"53",
         11144 => x"16",
         11145 => x"98",
         11146 => x"5c",
         11147 => x"94",
         11148 => x"8c",
         11149 => x"26",
         11150 => x"16",
         11151 => x"81",
         11152 => x"7c",
         11153 => x"94",
         11154 => x"56",
         11155 => x"1c",
         11156 => x"f8",
         11157 => x"08",
         11158 => x"ff",
         11159 => x"84",
         11160 => x"55",
         11161 => x"08",
         11162 => x"90",
         11163 => x"fd",
         11164 => x"52",
         11165 => x"ab",
         11166 => x"b8",
         11167 => x"84",
         11168 => x"fb",
         11169 => x"39",
         11170 => x"16",
         11171 => x"16",
         11172 => x"17",
         11173 => x"ff",
         11174 => x"84",
         11175 => x"81",
         11176 => x"b8",
         11177 => x"17",
         11178 => x"08",
         11179 => x"31",
         11180 => x"17",
         11181 => x"89",
         11182 => x"33",
         11183 => x"2e",
         11184 => x"fc",
         11185 => x"54",
         11186 => x"a0",
         11187 => x"53",
         11188 => x"16",
         11189 => x"96",
         11190 => x"56",
         11191 => x"81",
         11192 => x"ff",
         11193 => x"84",
         11194 => x"81",
         11195 => x"f9",
         11196 => x"7a",
         11197 => x"f9",
         11198 => x"54",
         11199 => x"53",
         11200 => x"53",
         11201 => x"52",
         11202 => x"c6",
         11203 => x"e4",
         11204 => x"38",
         11205 => x"08",
         11206 => x"b4",
         11207 => x"17",
         11208 => x"74",
         11209 => x"27",
         11210 => x"82",
         11211 => x"77",
         11212 => x"81",
         11213 => x"38",
         11214 => x"16",
         11215 => x"08",
         11216 => x"52",
         11217 => x"51",
         11218 => x"3f",
         11219 => x"12",
         11220 => x"08",
         11221 => x"f4",
         11222 => x"91",
         11223 => x"0b",
         11224 => x"0c",
         11225 => x"04",
         11226 => x"1b",
         11227 => x"84",
         11228 => x"92",
         11229 => x"f5",
         11230 => x"58",
         11231 => x"80",
         11232 => x"77",
         11233 => x"80",
         11234 => x"75",
         11235 => x"80",
         11236 => x"86",
         11237 => x"19",
         11238 => x"78",
         11239 => x"b5",
         11240 => x"74",
         11241 => x"79",
         11242 => x"90",
         11243 => x"86",
         11244 => x"5c",
         11245 => x"2e",
         11246 => x"7b",
         11247 => x"5a",
         11248 => x"08",
         11249 => x"38",
         11250 => x"5b",
         11251 => x"38",
         11252 => x"53",
         11253 => x"81",
         11254 => x"ff",
         11255 => x"84",
         11256 => x"80",
         11257 => x"ff",
         11258 => x"78",
         11259 => x"75",
         11260 => x"a4",
         11261 => x"11",
         11262 => x"5a",
         11263 => x"18",
         11264 => x"88",
         11265 => x"83",
         11266 => x"5d",
         11267 => x"9a",
         11268 => x"88",
         11269 => x"9b",
         11270 => x"17",
         11271 => x"19",
         11272 => x"74",
         11273 => x"c1",
         11274 => x"08",
         11275 => x"34",
         11276 => x"5b",
         11277 => x"34",
         11278 => x"56",
         11279 => x"34",
         11280 => x"59",
         11281 => x"34",
         11282 => x"80",
         11283 => x"34",
         11284 => x"18",
         11285 => x"0b",
         11286 => x"80",
         11287 => x"34",
         11288 => x"18",
         11289 => x"81",
         11290 => x"34",
         11291 => x"96",
         11292 => x"b8",
         11293 => x"19",
         11294 => x"06",
         11295 => x"90",
         11296 => x"84",
         11297 => x"8d",
         11298 => x"81",
         11299 => x"08",
         11300 => x"70",
         11301 => x"33",
         11302 => x"93",
         11303 => x"56",
         11304 => x"08",
         11305 => x"84",
         11306 => x"83",
         11307 => x"17",
         11308 => x"08",
         11309 => x"e4",
         11310 => x"74",
         11311 => x"27",
         11312 => x"82",
         11313 => x"74",
         11314 => x"81",
         11315 => x"38",
         11316 => x"17",
         11317 => x"08",
         11318 => x"52",
         11319 => x"51",
         11320 => x"3f",
         11321 => x"e8",
         11322 => x"2a",
         11323 => x"18",
         11324 => x"2a",
         11325 => x"18",
         11326 => x"08",
         11327 => x"34",
         11328 => x"5b",
         11329 => x"34",
         11330 => x"56",
         11331 => x"34",
         11332 => x"59",
         11333 => x"34",
         11334 => x"80",
         11335 => x"34",
         11336 => x"18",
         11337 => x"0b",
         11338 => x"80",
         11339 => x"34",
         11340 => x"18",
         11341 => x"81",
         11342 => x"34",
         11343 => x"94",
         11344 => x"b8",
         11345 => x"19",
         11346 => x"06",
         11347 => x"90",
         11348 => x"ae",
         11349 => x"33",
         11350 => x"a5",
         11351 => x"e4",
         11352 => x"55",
         11353 => x"38",
         11354 => x"56",
         11355 => x"39",
         11356 => x"79",
         11357 => x"fb",
         11358 => x"b8",
         11359 => x"84",
         11360 => x"b1",
         11361 => x"74",
         11362 => x"38",
         11363 => x"72",
         11364 => x"38",
         11365 => x"71",
         11366 => x"38",
         11367 => x"84",
         11368 => x"52",
         11369 => x"96",
         11370 => x"71",
         11371 => x"75",
         11372 => x"75",
         11373 => x"b8",
         11374 => x"3d",
         11375 => x"13",
         11376 => x"8f",
         11377 => x"b8",
         11378 => x"06",
         11379 => x"38",
         11380 => x"53",
         11381 => x"f6",
         11382 => x"7d",
         11383 => x"5b",
         11384 => x"b2",
         11385 => x"81",
         11386 => x"70",
         11387 => x"52",
         11388 => x"ac",
         11389 => x"38",
         11390 => x"a4",
         11391 => x"c0",
         11392 => x"71",
         11393 => x"70",
         11394 => x"34",
         11395 => x"b8",
         11396 => x"3d",
         11397 => x"0b",
         11398 => x"0c",
         11399 => x"04",
         11400 => x"11",
         11401 => x"06",
         11402 => x"70",
         11403 => x"38",
         11404 => x"81",
         11405 => x"05",
         11406 => x"76",
         11407 => x"38",
         11408 => x"e4",
         11409 => x"79",
         11410 => x"57",
         11411 => x"05",
         11412 => x"70",
         11413 => x"33",
         11414 => x"53",
         11415 => x"99",
         11416 => x"e0",
         11417 => x"ff",
         11418 => x"ff",
         11419 => x"70",
         11420 => x"38",
         11421 => x"81",
         11422 => x"54",
         11423 => x"9f",
         11424 => x"71",
         11425 => x"81",
         11426 => x"73",
         11427 => x"74",
         11428 => x"30",
         11429 => x"9f",
         11430 => x"59",
         11431 => x"80",
         11432 => x"81",
         11433 => x"5b",
         11434 => x"25",
         11435 => x"7a",
         11436 => x"39",
         11437 => x"f7",
         11438 => x"5e",
         11439 => x"39",
         11440 => x"80",
         11441 => x"cc",
         11442 => x"3d",
         11443 => x"3f",
         11444 => x"08",
         11445 => x"e4",
         11446 => x"8a",
         11447 => x"b8",
         11448 => x"3d",
         11449 => x"5c",
         11450 => x"3d",
         11451 => x"c5",
         11452 => x"b8",
         11453 => x"84",
         11454 => x"80",
         11455 => x"80",
         11456 => x"70",
         11457 => x"5a",
         11458 => x"80",
         11459 => x"b2",
         11460 => x"84",
         11461 => x"57",
         11462 => x"2e",
         11463 => x"63",
         11464 => x"9a",
         11465 => x"88",
         11466 => x"33",
         11467 => x"57",
         11468 => x"2e",
         11469 => x"98",
         11470 => x"84",
         11471 => x"98",
         11472 => x"84",
         11473 => x"84",
         11474 => x"06",
         11475 => x"85",
         11476 => x"e4",
         11477 => x"0d",
         11478 => x"33",
         11479 => x"71",
         11480 => x"90",
         11481 => x"07",
         11482 => x"5b",
         11483 => x"7a",
         11484 => x"0c",
         11485 => x"b8",
         11486 => x"3d",
         11487 => x"9e",
         11488 => x"e6",
         11489 => x"e6",
         11490 => x"40",
         11491 => x"80",
         11492 => x"3d",
         11493 => x"52",
         11494 => x"51",
         11495 => x"84",
         11496 => x"59",
         11497 => x"08",
         11498 => x"60",
         11499 => x"0c",
         11500 => x"11",
         11501 => x"3d",
         11502 => x"db",
         11503 => x"58",
         11504 => x"82",
         11505 => x"d8",
         11506 => x"40",
         11507 => x"7a",
         11508 => x"aa",
         11509 => x"e4",
         11510 => x"b8",
         11511 => x"92",
         11512 => x"df",
         11513 => x"56",
         11514 => x"77",
         11515 => x"84",
         11516 => x"83",
         11517 => x"5d",
         11518 => x"38",
         11519 => x"53",
         11520 => x"81",
         11521 => x"ff",
         11522 => x"84",
         11523 => x"80",
         11524 => x"ff",
         11525 => x"76",
         11526 => x"78",
         11527 => x"80",
         11528 => x"9b",
         11529 => x"12",
         11530 => x"2b",
         11531 => x"33",
         11532 => x"56",
         11533 => x"2e",
         11534 => x"76",
         11535 => x"0c",
         11536 => x"51",
         11537 => x"3f",
         11538 => x"08",
         11539 => x"e4",
         11540 => x"38",
         11541 => x"51",
         11542 => x"3f",
         11543 => x"08",
         11544 => x"e4",
         11545 => x"80",
         11546 => x"9b",
         11547 => x"12",
         11548 => x"2b",
         11549 => x"33",
         11550 => x"5e",
         11551 => x"2e",
         11552 => x"76",
         11553 => x"38",
         11554 => x"08",
         11555 => x"ff",
         11556 => x"84",
         11557 => x"59",
         11558 => x"08",
         11559 => x"b4",
         11560 => x"2e",
         11561 => x"78",
         11562 => x"80",
         11563 => x"b8",
         11564 => x"51",
         11565 => x"3f",
         11566 => x"05",
         11567 => x"79",
         11568 => x"38",
         11569 => x"81",
         11570 => x"70",
         11571 => x"57",
         11572 => x"81",
         11573 => x"78",
         11574 => x"38",
         11575 => x"9c",
         11576 => x"82",
         11577 => x"18",
         11578 => x"08",
         11579 => x"ff",
         11580 => x"56",
         11581 => x"75",
         11582 => x"38",
         11583 => x"e6",
         11584 => x"5f",
         11585 => x"34",
         11586 => x"08",
         11587 => x"bd",
         11588 => x"2e",
         11589 => x"80",
         11590 => x"c0",
         11591 => x"10",
         11592 => x"05",
         11593 => x"33",
         11594 => x"5e",
         11595 => x"2e",
         11596 => x"1a",
         11597 => x"33",
         11598 => x"74",
         11599 => x"1a",
         11600 => x"26",
         11601 => x"57",
         11602 => x"94",
         11603 => x"5f",
         11604 => x"70",
         11605 => x"34",
         11606 => x"79",
         11607 => x"38",
         11608 => x"81",
         11609 => x"76",
         11610 => x"81",
         11611 => x"38",
         11612 => x"7c",
         11613 => x"b8",
         11614 => x"e4",
         11615 => x"95",
         11616 => x"17",
         11617 => x"2b",
         11618 => x"07",
         11619 => x"56",
         11620 => x"39",
         11621 => x"94",
         11622 => x"98",
         11623 => x"2b",
         11624 => x"80",
         11625 => x"5a",
         11626 => x"7a",
         11627 => x"ce",
         11628 => x"e4",
         11629 => x"b8",
         11630 => x"2e",
         11631 => x"ff",
         11632 => x"54",
         11633 => x"53",
         11634 => x"53",
         11635 => x"52",
         11636 => x"fe",
         11637 => x"84",
         11638 => x"fc",
         11639 => x"b8",
         11640 => x"17",
         11641 => x"08",
         11642 => x"31",
         11643 => x"08",
         11644 => x"a0",
         11645 => x"fc",
         11646 => x"16",
         11647 => x"82",
         11648 => x"06",
         11649 => x"81",
         11650 => x"08",
         11651 => x"05",
         11652 => x"81",
         11653 => x"ff",
         11654 => x"7c",
         11655 => x"39",
         11656 => x"e6",
         11657 => x"5c",
         11658 => x"34",
         11659 => x"d0",
         11660 => x"10",
         11661 => x"d4",
         11662 => x"70",
         11663 => x"59",
         11664 => x"7a",
         11665 => x"06",
         11666 => x"fd",
         11667 => x"e5",
         11668 => x"81",
         11669 => x"79",
         11670 => x"81",
         11671 => x"77",
         11672 => x"8e",
         11673 => x"3d",
         11674 => x"19",
         11675 => x"33",
         11676 => x"05",
         11677 => x"78",
         11678 => x"fd",
         11679 => x"59",
         11680 => x"78",
         11681 => x"0c",
         11682 => x"0d",
         11683 => x"0d",
         11684 => x"55",
         11685 => x"80",
         11686 => x"74",
         11687 => x"80",
         11688 => x"73",
         11689 => x"80",
         11690 => x"86",
         11691 => x"16",
         11692 => x"78",
         11693 => x"a0",
         11694 => x"72",
         11695 => x"75",
         11696 => x"91",
         11697 => x"72",
         11698 => x"8c",
         11699 => x"76",
         11700 => x"b9",
         11701 => x"08",
         11702 => x"76",
         11703 => x"cc",
         11704 => x"11",
         11705 => x"2b",
         11706 => x"73",
         11707 => x"f7",
         11708 => x"ff",
         11709 => x"bb",
         11710 => x"b8",
         11711 => x"15",
         11712 => x"53",
         11713 => x"bb",
         11714 => x"b8",
         11715 => x"26",
         11716 => x"75",
         11717 => x"70",
         11718 => x"77",
         11719 => x"17",
         11720 => x"59",
         11721 => x"82",
         11722 => x"77",
         11723 => x"38",
         11724 => x"94",
         11725 => x"94",
         11726 => x"16",
         11727 => x"2a",
         11728 => x"5a",
         11729 => x"2e",
         11730 => x"73",
         11731 => x"ff",
         11732 => x"84",
         11733 => x"54",
         11734 => x"08",
         11735 => x"a3",
         11736 => x"2e",
         11737 => x"74",
         11738 => x"38",
         11739 => x"9c",
         11740 => x"82",
         11741 => x"98",
         11742 => x"ae",
         11743 => x"91",
         11744 => x"53",
         11745 => x"e4",
         11746 => x"0d",
         11747 => x"33",
         11748 => x"81",
         11749 => x"73",
         11750 => x"75",
         11751 => x"55",
         11752 => x"76",
         11753 => x"81",
         11754 => x"38",
         11755 => x"0c",
         11756 => x"54",
         11757 => x"90",
         11758 => x"16",
         11759 => x"33",
         11760 => x"57",
         11761 => x"34",
         11762 => x"06",
         11763 => x"2e",
         11764 => x"15",
         11765 => x"85",
         11766 => x"16",
         11767 => x"84",
         11768 => x"8b",
         11769 => x"80",
         11770 => x"0c",
         11771 => x"54",
         11772 => x"80",
         11773 => x"98",
         11774 => x"80",
         11775 => x"38",
         11776 => x"84",
         11777 => x"57",
         11778 => x"17",
         11779 => x"76",
         11780 => x"56",
         11781 => x"a9",
         11782 => x"15",
         11783 => x"fe",
         11784 => x"56",
         11785 => x"80",
         11786 => x"16",
         11787 => x"29",
         11788 => x"05",
         11789 => x"11",
         11790 => x"78",
         11791 => x"df",
         11792 => x"08",
         11793 => x"39",
         11794 => x"51",
         11795 => x"3f",
         11796 => x"08",
         11797 => x"39",
         11798 => x"51",
         11799 => x"3f",
         11800 => x"08",
         11801 => x"72",
         11802 => x"72",
         11803 => x"56",
         11804 => x"73",
         11805 => x"ff",
         11806 => x"84",
         11807 => x"54",
         11808 => x"08",
         11809 => x"38",
         11810 => x"08",
         11811 => x"ed",
         11812 => x"e4",
         11813 => x"0c",
         11814 => x"0c",
         11815 => x"82",
         11816 => x"34",
         11817 => x"b8",
         11818 => x"3d",
         11819 => x"3d",
         11820 => x"89",
         11821 => x"2e",
         11822 => x"53",
         11823 => x"05",
         11824 => x"84",
         11825 => x"9b",
         11826 => x"e4",
         11827 => x"b8",
         11828 => x"2e",
         11829 => x"76",
         11830 => x"73",
         11831 => x"0c",
         11832 => x"04",
         11833 => x"7d",
         11834 => x"ff",
         11835 => x"84",
         11836 => x"55",
         11837 => x"08",
         11838 => x"ab",
         11839 => x"98",
         11840 => x"80",
         11841 => x"38",
         11842 => x"70",
         11843 => x"06",
         11844 => x"80",
         11845 => x"38",
         11846 => x"9b",
         11847 => x"12",
         11848 => x"2b",
         11849 => x"33",
         11850 => x"55",
         11851 => x"2e",
         11852 => x"88",
         11853 => x"58",
         11854 => x"84",
         11855 => x"52",
         11856 => x"99",
         11857 => x"b8",
         11858 => x"74",
         11859 => x"38",
         11860 => x"ff",
         11861 => x"76",
         11862 => x"39",
         11863 => x"76",
         11864 => x"39",
         11865 => x"94",
         11866 => x"98",
         11867 => x"2b",
         11868 => x"88",
         11869 => x"5a",
         11870 => x"fa",
         11871 => x"55",
         11872 => x"80",
         11873 => x"74",
         11874 => x"80",
         11875 => x"72",
         11876 => x"80",
         11877 => x"86",
         11878 => x"16",
         11879 => x"71",
         11880 => x"38",
         11881 => x"57",
         11882 => x"73",
         11883 => x"84",
         11884 => x"88",
         11885 => x"81",
         11886 => x"fe",
         11887 => x"84",
         11888 => x"81",
         11889 => x"dc",
         11890 => x"08",
         11891 => x"39",
         11892 => x"7a",
         11893 => x"89",
         11894 => x"2e",
         11895 => x"08",
         11896 => x"2e",
         11897 => x"33",
         11898 => x"2e",
         11899 => x"14",
         11900 => x"22",
         11901 => x"78",
         11902 => x"38",
         11903 => x"59",
         11904 => x"80",
         11905 => x"80",
         11906 => x"38",
         11907 => x"51",
         11908 => x"3f",
         11909 => x"08",
         11910 => x"e4",
         11911 => x"b5",
         11912 => x"e4",
         11913 => x"76",
         11914 => x"ff",
         11915 => x"72",
         11916 => x"ff",
         11917 => x"84",
         11918 => x"84",
         11919 => x"70",
         11920 => x"2c",
         11921 => x"08",
         11922 => x"54",
         11923 => x"e4",
         11924 => x"0d",
         11925 => x"53",
         11926 => x"ff",
         11927 => x"72",
         11928 => x"ff",
         11929 => x"84",
         11930 => x"84",
         11931 => x"70",
         11932 => x"2c",
         11933 => x"08",
         11934 => x"54",
         11935 => x"52",
         11936 => x"96",
         11937 => x"b8",
         11938 => x"b8",
         11939 => x"3d",
         11940 => x"14",
         11941 => x"fd",
         11942 => x"b8",
         11943 => x"06",
         11944 => x"d8",
         11945 => x"08",
         11946 => x"d2",
         11947 => x"0d",
         11948 => x"53",
         11949 => x"53",
         11950 => x"56",
         11951 => x"84",
         11952 => x"55",
         11953 => x"08",
         11954 => x"38",
         11955 => x"e4",
         11956 => x"0d",
         11957 => x"75",
         11958 => x"a9",
         11959 => x"e4",
         11960 => x"b8",
         11961 => x"38",
         11962 => x"05",
         11963 => x"2b",
         11964 => x"74",
         11965 => x"76",
         11966 => x"38",
         11967 => x"51",
         11968 => x"3f",
         11969 => x"e4",
         11970 => x"0d",
         11971 => x"84",
         11972 => x"95",
         11973 => x"ed",
         11974 => x"68",
         11975 => x"53",
         11976 => x"05",
         11977 => x"51",
         11978 => x"84",
         11979 => x"5a",
         11980 => x"08",
         11981 => x"75",
         11982 => x"9c",
         11983 => x"11",
         11984 => x"59",
         11985 => x"75",
         11986 => x"38",
         11987 => x"79",
         11988 => x"0c",
         11989 => x"04",
         11990 => x"08",
         11991 => x"5b",
         11992 => x"82",
         11993 => x"a8",
         11994 => x"b8",
         11995 => x"5d",
         11996 => x"c1",
         11997 => x"1d",
         11998 => x"56",
         11999 => x"76",
         12000 => x"38",
         12001 => x"78",
         12002 => x"81",
         12003 => x"54",
         12004 => x"17",
         12005 => x"33",
         12006 => x"b7",
         12007 => x"e4",
         12008 => x"85",
         12009 => x"81",
         12010 => x"18",
         12011 => x"5b",
         12012 => x"cc",
         12013 => x"5e",
         12014 => x"82",
         12015 => x"17",
         12016 => x"11",
         12017 => x"33",
         12018 => x"71",
         12019 => x"81",
         12020 => x"72",
         12021 => x"75",
         12022 => x"ff",
         12023 => x"06",
         12024 => x"70",
         12025 => x"05",
         12026 => x"83",
         12027 => x"ff",
         12028 => x"43",
         12029 => x"53",
         12030 => x"56",
         12031 => x"38",
         12032 => x"7a",
         12033 => x"84",
         12034 => x"07",
         12035 => x"18",
         12036 => x"b8",
         12037 => x"3d",
         12038 => x"54",
         12039 => x"53",
         12040 => x"53",
         12041 => x"52",
         12042 => x"a6",
         12043 => x"84",
         12044 => x"fe",
         12045 => x"b8",
         12046 => x"18",
         12047 => x"08",
         12048 => x"31",
         12049 => x"08",
         12050 => x"a0",
         12051 => x"fe",
         12052 => x"17",
         12053 => x"82",
         12054 => x"06",
         12055 => x"81",
         12056 => x"08",
         12057 => x"05",
         12058 => x"81",
         12059 => x"fe",
         12060 => x"77",
         12061 => x"39",
         12062 => x"92",
         12063 => x"75",
         12064 => x"ff",
         12065 => x"84",
         12066 => x"ff",
         12067 => x"38",
         12068 => x"08",
         12069 => x"f7",
         12070 => x"e4",
         12071 => x"84",
         12072 => x"07",
         12073 => x"05",
         12074 => x"5a",
         12075 => x"9c",
         12076 => x"26",
         12077 => x"7f",
         12078 => x"18",
         12079 => x"33",
         12080 => x"77",
         12081 => x"fe",
         12082 => x"17",
         12083 => x"11",
         12084 => x"71",
         12085 => x"70",
         12086 => x"25",
         12087 => x"83",
         12088 => x"1f",
         12089 => x"59",
         12090 => x"78",
         12091 => x"fe",
         12092 => x"5a",
         12093 => x"81",
         12094 => x"7a",
         12095 => x"94",
         12096 => x"17",
         12097 => x"58",
         12098 => x"34",
         12099 => x"82",
         12100 => x"e7",
         12101 => x"0d",
         12102 => x"56",
         12103 => x"9f",
         12104 => x"55",
         12105 => x"97",
         12106 => x"54",
         12107 => x"8f",
         12108 => x"22",
         12109 => x"59",
         12110 => x"2e",
         12111 => x"80",
         12112 => x"75",
         12113 => x"91",
         12114 => x"75",
         12115 => x"90",
         12116 => x"81",
         12117 => x"55",
         12118 => x"73",
         12119 => x"c4",
         12120 => x"08",
         12121 => x"18",
         12122 => x"38",
         12123 => x"38",
         12124 => x"77",
         12125 => x"81",
         12126 => x"38",
         12127 => x"74",
         12128 => x"82",
         12129 => x"88",
         12130 => x"17",
         12131 => x"0c",
         12132 => x"07",
         12133 => x"18",
         12134 => x"2e",
         12135 => x"91",
         12136 => x"55",
         12137 => x"e4",
         12138 => x"0d",
         12139 => x"78",
         12140 => x"ff",
         12141 => x"76",
         12142 => x"ca",
         12143 => x"e4",
         12144 => x"b8",
         12145 => x"2e",
         12146 => x"84",
         12147 => x"81",
         12148 => x"38",
         12149 => x"08",
         12150 => x"e5",
         12151 => x"73",
         12152 => x"ff",
         12153 => x"84",
         12154 => x"82",
         12155 => x"16",
         12156 => x"94",
         12157 => x"55",
         12158 => x"27",
         12159 => x"81",
         12160 => x"0c",
         12161 => x"81",
         12162 => x"84",
         12163 => x"54",
         12164 => x"ff",
         12165 => x"39",
         12166 => x"51",
         12167 => x"3f",
         12168 => x"08",
         12169 => x"73",
         12170 => x"73",
         12171 => x"56",
         12172 => x"80",
         12173 => x"33",
         12174 => x"56",
         12175 => x"18",
         12176 => x"39",
         12177 => x"52",
         12178 => x"fd",
         12179 => x"b8",
         12180 => x"2e",
         12181 => x"84",
         12182 => x"81",
         12183 => x"38",
         12184 => x"38",
         12185 => x"b8",
         12186 => x"19",
         12187 => x"a1",
         12188 => x"e4",
         12189 => x"08",
         12190 => x"56",
         12191 => x"84",
         12192 => x"27",
         12193 => x"84",
         12194 => x"9c",
         12195 => x"81",
         12196 => x"80",
         12197 => x"ff",
         12198 => x"75",
         12199 => x"c7",
         12200 => x"e4",
         12201 => x"b8",
         12202 => x"e3",
         12203 => x"76",
         12204 => x"d2",
         12205 => x"e4",
         12206 => x"b8",
         12207 => x"2e",
         12208 => x"84",
         12209 => x"81",
         12210 => x"38",
         12211 => x"08",
         12212 => x"fe",
         12213 => x"73",
         12214 => x"ff",
         12215 => x"84",
         12216 => x"80",
         12217 => x"16",
         12218 => x"94",
         12219 => x"55",
         12220 => x"27",
         12221 => x"15",
         12222 => x"84",
         12223 => x"07",
         12224 => x"17",
         12225 => x"77",
         12226 => x"a1",
         12227 => x"74",
         12228 => x"33",
         12229 => x"39",
         12230 => x"bb",
         12231 => x"90",
         12232 => x"56",
         12233 => x"82",
         12234 => x"82",
         12235 => x"33",
         12236 => x"86",
         12237 => x"e4",
         12238 => x"33",
         12239 => x"fa",
         12240 => x"90",
         12241 => x"54",
         12242 => x"84",
         12243 => x"56",
         12244 => x"56",
         12245 => x"db",
         12246 => x"53",
         12247 => x"9c",
         12248 => x"3d",
         12249 => x"fb",
         12250 => x"e4",
         12251 => x"b8",
         12252 => x"2e",
         12253 => x"84",
         12254 => x"a7",
         12255 => x"7d",
         12256 => x"08",
         12257 => x"70",
         12258 => x"ab",
         12259 => x"b8",
         12260 => x"84",
         12261 => x"de",
         12262 => x"93",
         12263 => x"85",
         12264 => x"59",
         12265 => x"77",
         12266 => x"98",
         12267 => x"7b",
         12268 => x"02",
         12269 => x"33",
         12270 => x"5d",
         12271 => x"7b",
         12272 => x"7d",
         12273 => x"9b",
         12274 => x"12",
         12275 => x"2b",
         12276 => x"41",
         12277 => x"58",
         12278 => x"80",
         12279 => x"84",
         12280 => x"57",
         12281 => x"80",
         12282 => x"56",
         12283 => x"7b",
         12284 => x"38",
         12285 => x"41",
         12286 => x"08",
         12287 => x"70",
         12288 => x"8b",
         12289 => x"b8",
         12290 => x"84",
         12291 => x"fe",
         12292 => x"b8",
         12293 => x"74",
         12294 => x"b4",
         12295 => x"e4",
         12296 => x"b8",
         12297 => x"38",
         12298 => x"b8",
         12299 => x"3d",
         12300 => x"16",
         12301 => x"33",
         12302 => x"71",
         12303 => x"7d",
         12304 => x"5d",
         12305 => x"84",
         12306 => x"84",
         12307 => x"84",
         12308 => x"fe",
         12309 => x"08",
         12310 => x"08",
         12311 => x"74",
         12312 => x"d3",
         12313 => x"78",
         12314 => x"92",
         12315 => x"e4",
         12316 => x"b8",
         12317 => x"2e",
         12318 => x"30",
         12319 => x"80",
         12320 => x"7a",
         12321 => x"38",
         12322 => x"95",
         12323 => x"08",
         12324 => x"7b",
         12325 => x"9c",
         12326 => x"26",
         12327 => x"82",
         12328 => x"d2",
         12329 => x"fe",
         12330 => x"84",
         12331 => x"84",
         12332 => x"a7",
         12333 => x"b8",
         12334 => x"19",
         12335 => x"5a",
         12336 => x"76",
         12337 => x"38",
         12338 => x"7a",
         12339 => x"7a",
         12340 => x"06",
         12341 => x"81",
         12342 => x"b8",
         12343 => x"17",
         12344 => x"f1",
         12345 => x"b8",
         12346 => x"2e",
         12347 => x"56",
         12348 => x"b4",
         12349 => x"56",
         12350 => x"9c",
         12351 => x"e5",
         12352 => x"0b",
         12353 => x"90",
         12354 => x"27",
         12355 => x"80",
         12356 => x"ff",
         12357 => x"84",
         12358 => x"56",
         12359 => x"08",
         12360 => x"96",
         12361 => x"2e",
         12362 => x"fe",
         12363 => x"56",
         12364 => x"81",
         12365 => x"08",
         12366 => x"81",
         12367 => x"fe",
         12368 => x"81",
         12369 => x"e4",
         12370 => x"09",
         12371 => x"a6",
         12372 => x"e4",
         12373 => x"34",
         12374 => x"a8",
         12375 => x"84",
         12376 => x"59",
         12377 => x"18",
         12378 => x"eb",
         12379 => x"33",
         12380 => x"2e",
         12381 => x"fe",
         12382 => x"54",
         12383 => x"a0",
         12384 => x"53",
         12385 => x"17",
         12386 => x"f1",
         12387 => x"58",
         12388 => x"79",
         12389 => x"27",
         12390 => x"74",
         12391 => x"fe",
         12392 => x"84",
         12393 => x"5a",
         12394 => x"08",
         12395 => x"cb",
         12396 => x"e4",
         12397 => x"fd",
         12398 => x"b8",
         12399 => x"2e",
         12400 => x"80",
         12401 => x"76",
         12402 => x"9b",
         12403 => x"e4",
         12404 => x"9c",
         12405 => x"11",
         12406 => x"58",
         12407 => x"7b",
         12408 => x"38",
         12409 => x"18",
         12410 => x"33",
         12411 => x"7b",
         12412 => x"79",
         12413 => x"26",
         12414 => x"80",
         12415 => x"39",
         12416 => x"f7",
         12417 => x"e4",
         12418 => x"95",
         12419 => x"fd",
         12420 => x"3d",
         12421 => x"9f",
         12422 => x"05",
         12423 => x"51",
         12424 => x"3f",
         12425 => x"08",
         12426 => x"e4",
         12427 => x"8a",
         12428 => x"b8",
         12429 => x"3d",
         12430 => x"43",
         12431 => x"3d",
         12432 => x"ff",
         12433 => x"84",
         12434 => x"56",
         12435 => x"08",
         12436 => x"0b",
         12437 => x"0c",
         12438 => x"04",
         12439 => x"08",
         12440 => x"81",
         12441 => x"02",
         12442 => x"33",
         12443 => x"81",
         12444 => x"86",
         12445 => x"b9",
         12446 => x"74",
         12447 => x"70",
         12448 => x"83",
         12449 => x"b8",
         12450 => x"57",
         12451 => x"e4",
         12452 => x"87",
         12453 => x"e4",
         12454 => x"80",
         12455 => x"b8",
         12456 => x"2e",
         12457 => x"75",
         12458 => x"7d",
         12459 => x"08",
         12460 => x"5d",
         12461 => x"80",
         12462 => x"19",
         12463 => x"fe",
         12464 => x"80",
         12465 => x"27",
         12466 => x"17",
         12467 => x"29",
         12468 => x"05",
         12469 => x"b4",
         12470 => x"17",
         12471 => x"79",
         12472 => x"76",
         12473 => x"58",
         12474 => x"55",
         12475 => x"74",
         12476 => x"22",
         12477 => x"27",
         12478 => x"81",
         12479 => x"53",
         12480 => x"17",
         12481 => x"ee",
         12482 => x"b8",
         12483 => x"df",
         12484 => x"58",
         12485 => x"56",
         12486 => x"81",
         12487 => x"08",
         12488 => x"70",
         12489 => x"33",
         12490 => x"ee",
         12491 => x"56",
         12492 => x"08",
         12493 => x"b8",
         12494 => x"18",
         12495 => x"08",
         12496 => x"31",
         12497 => x"18",
         12498 => x"ee",
         12499 => x"33",
         12500 => x"2e",
         12501 => x"fe",
         12502 => x"54",
         12503 => x"a0",
         12504 => x"53",
         12505 => x"17",
         12506 => x"ed",
         12507 => x"ca",
         12508 => x"7b",
         12509 => x"55",
         12510 => x"fd",
         12511 => x"9c",
         12512 => x"fd",
         12513 => x"52",
         12514 => x"f2",
         12515 => x"b8",
         12516 => x"84",
         12517 => x"80",
         12518 => x"38",
         12519 => x"08",
         12520 => x"8d",
         12521 => x"e4",
         12522 => x"fd",
         12523 => x"53",
         12524 => x"51",
         12525 => x"3f",
         12526 => x"08",
         12527 => x"9c",
         12528 => x"11",
         12529 => x"5a",
         12530 => x"7b",
         12531 => x"81",
         12532 => x"0c",
         12533 => x"81",
         12534 => x"84",
         12535 => x"55",
         12536 => x"ff",
         12537 => x"84",
         12538 => x"9f",
         12539 => x"8a",
         12540 => x"74",
         12541 => x"06",
         12542 => x"76",
         12543 => x"81",
         12544 => x"38",
         12545 => x"1f",
         12546 => x"75",
         12547 => x"57",
         12548 => x"56",
         12549 => x"7d",
         12550 => x"b8",
         12551 => x"58",
         12552 => x"c3",
         12553 => x"59",
         12554 => x"1a",
         12555 => x"cf",
         12556 => x"0b",
         12557 => x"34",
         12558 => x"80",
         12559 => x"7d",
         12560 => x"ff",
         12561 => x"77",
         12562 => x"34",
         12563 => x"5b",
         12564 => x"17",
         12565 => x"55",
         12566 => x"81",
         12567 => x"59",
         12568 => x"d8",
         12569 => x"57",
         12570 => x"70",
         12571 => x"33",
         12572 => x"05",
         12573 => x"16",
         12574 => x"38",
         12575 => x"0b",
         12576 => x"34",
         12577 => x"83",
         12578 => x"5b",
         12579 => x"80",
         12580 => x"78",
         12581 => x"7a",
         12582 => x"34",
         12583 => x"74",
         12584 => x"f0",
         12585 => x"81",
         12586 => x"34",
         12587 => x"92",
         12588 => x"b8",
         12589 => x"84",
         12590 => x"fd",
         12591 => x"56",
         12592 => x"08",
         12593 => x"84",
         12594 => x"97",
         12595 => x"0b",
         12596 => x"80",
         12597 => x"17",
         12598 => x"58",
         12599 => x"18",
         12600 => x"2a",
         12601 => x"18",
         12602 => x"5a",
         12603 => x"80",
         12604 => x"55",
         12605 => x"16",
         12606 => x"81",
         12607 => x"34",
         12608 => x"ed",
         12609 => x"b8",
         12610 => x"75",
         12611 => x"0c",
         12612 => x"04",
         12613 => x"55",
         12614 => x"17",
         12615 => x"2a",
         12616 => x"ed",
         12617 => x"fd",
         12618 => x"2a",
         12619 => x"cc",
         12620 => x"88",
         12621 => x"80",
         12622 => x"7d",
         12623 => x"80",
         12624 => x"1b",
         12625 => x"fe",
         12626 => x"90",
         12627 => x"94",
         12628 => x"88",
         12629 => x"95",
         12630 => x"55",
         12631 => x"16",
         12632 => x"81",
         12633 => x"34",
         12634 => x"ec",
         12635 => x"b8",
         12636 => x"ff",
         12637 => x"3d",
         12638 => x"b4",
         12639 => x"59",
         12640 => x"80",
         12641 => x"79",
         12642 => x"5b",
         12643 => x"26",
         12644 => x"ba",
         12645 => x"38",
         12646 => x"75",
         12647 => x"af",
         12648 => x"b1",
         12649 => x"05",
         12650 => x"51",
         12651 => x"3f",
         12652 => x"08",
         12653 => x"e4",
         12654 => x"8a",
         12655 => x"b8",
         12656 => x"3d",
         12657 => x"a6",
         12658 => x"3d",
         12659 => x"3d",
         12660 => x"ff",
         12661 => x"84",
         12662 => x"56",
         12663 => x"08",
         12664 => x"81",
         12665 => x"81",
         12666 => x"86",
         12667 => x"38",
         12668 => x"3d",
         12669 => x"58",
         12670 => x"70",
         12671 => x"33",
         12672 => x"05",
         12673 => x"15",
         12674 => x"38",
         12675 => x"b0",
         12676 => x"58",
         12677 => x"81",
         12678 => x"77",
         12679 => x"59",
         12680 => x"55",
         12681 => x"b3",
         12682 => x"77",
         12683 => x"d5",
         12684 => x"e4",
         12685 => x"b8",
         12686 => x"d8",
         12687 => x"3d",
         12688 => x"cb",
         12689 => x"84",
         12690 => x"b1",
         12691 => x"76",
         12692 => x"70",
         12693 => x"57",
         12694 => x"89",
         12695 => x"82",
         12696 => x"ff",
         12697 => x"5d",
         12698 => x"2e",
         12699 => x"80",
         12700 => x"e4",
         12701 => x"72",
         12702 => x"5f",
         12703 => x"81",
         12704 => x"79",
         12705 => x"5b",
         12706 => x"12",
         12707 => x"77",
         12708 => x"38",
         12709 => x"81",
         12710 => x"55",
         12711 => x"58",
         12712 => x"89",
         12713 => x"70",
         12714 => x"58",
         12715 => x"70",
         12716 => x"55",
         12717 => x"09",
         12718 => x"38",
         12719 => x"38",
         12720 => x"70",
         12721 => x"07",
         12722 => x"07",
         12723 => x"7a",
         12724 => x"38",
         12725 => x"1e",
         12726 => x"83",
         12727 => x"38",
         12728 => x"5a",
         12729 => x"39",
         12730 => x"fd",
         12731 => x"7f",
         12732 => x"b1",
         12733 => x"05",
         12734 => x"51",
         12735 => x"3f",
         12736 => x"08",
         12737 => x"e4",
         12738 => x"38",
         12739 => x"6c",
         12740 => x"2e",
         12741 => x"fe",
         12742 => x"51",
         12743 => x"3f",
         12744 => x"08",
         12745 => x"e4",
         12746 => x"38",
         12747 => x"0b",
         12748 => x"88",
         12749 => x"05",
         12750 => x"75",
         12751 => x"57",
         12752 => x"81",
         12753 => x"ff",
         12754 => x"ef",
         12755 => x"cb",
         12756 => x"19",
         12757 => x"33",
         12758 => x"81",
         12759 => x"7e",
         12760 => x"a0",
         12761 => x"8b",
         12762 => x"5d",
         12763 => x"1e",
         12764 => x"33",
         12765 => x"81",
         12766 => x"75",
         12767 => x"c5",
         12768 => x"08",
         12769 => x"bd",
         12770 => x"19",
         12771 => x"33",
         12772 => x"07",
         12773 => x"58",
         12774 => x"83",
         12775 => x"38",
         12776 => x"18",
         12777 => x"5e",
         12778 => x"27",
         12779 => x"8a",
         12780 => x"71",
         12781 => x"08",
         12782 => x"75",
         12783 => x"b5",
         12784 => x"5d",
         12785 => x"08",
         12786 => x"38",
         12787 => x"5f",
         12788 => x"38",
         12789 => x"53",
         12790 => x"81",
         12791 => x"fe",
         12792 => x"84",
         12793 => x"80",
         12794 => x"ff",
         12795 => x"77",
         12796 => x"7f",
         12797 => x"d8",
         12798 => x"7b",
         12799 => x"81",
         12800 => x"79",
         12801 => x"81",
         12802 => x"6a",
         12803 => x"ff",
         12804 => x"7b",
         12805 => x"34",
         12806 => x"58",
         12807 => x"18",
         12808 => x"5b",
         12809 => x"09",
         12810 => x"38",
         12811 => x"5e",
         12812 => x"18",
         12813 => x"2a",
         12814 => x"ed",
         12815 => x"57",
         12816 => x"18",
         12817 => x"aa",
         12818 => x"3d",
         12819 => x"56",
         12820 => x"95",
         12821 => x"78",
         12822 => x"a2",
         12823 => x"e4",
         12824 => x"b8",
         12825 => x"f5",
         12826 => x"5c",
         12827 => x"57",
         12828 => x"16",
         12829 => x"b4",
         12830 => x"33",
         12831 => x"7e",
         12832 => x"81",
         12833 => x"38",
         12834 => x"53",
         12835 => x"81",
         12836 => x"fe",
         12837 => x"84",
         12838 => x"80",
         12839 => x"ff",
         12840 => x"76",
         12841 => x"77",
         12842 => x"38",
         12843 => x"5a",
         12844 => x"81",
         12845 => x"34",
         12846 => x"7b",
         12847 => x"80",
         12848 => x"fe",
         12849 => x"84",
         12850 => x"55",
         12851 => x"08",
         12852 => x"98",
         12853 => x"74",
         12854 => x"e1",
         12855 => x"74",
         12856 => x"7f",
         12857 => x"9d",
         12858 => x"e4",
         12859 => x"e4",
         12860 => x"0d",
         12861 => x"84",
         12862 => x"b1",
         12863 => x"95",
         12864 => x"19",
         12865 => x"2b",
         12866 => x"07",
         12867 => x"56",
         12868 => x"39",
         12869 => x"08",
         12870 => x"fe",
         12871 => x"e4",
         12872 => x"fe",
         12873 => x"84",
         12874 => x"b1",
         12875 => x"81",
         12876 => x"08",
         12877 => x"81",
         12878 => x"fe",
         12879 => x"81",
         12880 => x"e4",
         12881 => x"09",
         12882 => x"db",
         12883 => x"e4",
         12884 => x"34",
         12885 => x"a8",
         12886 => x"84",
         12887 => x"59",
         12888 => x"17",
         12889 => x"a0",
         12890 => x"33",
         12891 => x"2e",
         12892 => x"fe",
         12893 => x"54",
         12894 => x"a0",
         12895 => x"53",
         12896 => x"16",
         12897 => x"e1",
         12898 => x"58",
         12899 => x"81",
         12900 => x"08",
         12901 => x"70",
         12902 => x"33",
         12903 => x"e1",
         12904 => x"5c",
         12905 => x"08",
         12906 => x"84",
         12907 => x"83",
         12908 => x"17",
         12909 => x"08",
         12910 => x"e4",
         12911 => x"74",
         12912 => x"27",
         12913 => x"82",
         12914 => x"7c",
         12915 => x"81",
         12916 => x"38",
         12917 => x"17",
         12918 => x"08",
         12919 => x"52",
         12920 => x"51",
         12921 => x"3f",
         12922 => x"e8",
         12923 => x"0d",
         12924 => x"05",
         12925 => x"05",
         12926 => x"33",
         12927 => x"53",
         12928 => x"05",
         12929 => x"51",
         12930 => x"3f",
         12931 => x"08",
         12932 => x"e4",
         12933 => x"8a",
         12934 => x"b8",
         12935 => x"3d",
         12936 => x"5a",
         12937 => x"3d",
         12938 => x"ff",
         12939 => x"84",
         12940 => x"56",
         12941 => x"08",
         12942 => x"80",
         12943 => x"81",
         12944 => x"86",
         12945 => x"38",
         12946 => x"61",
         12947 => x"12",
         12948 => x"7a",
         12949 => x"51",
         12950 => x"73",
         12951 => x"78",
         12952 => x"83",
         12953 => x"51",
         12954 => x"3f",
         12955 => x"08",
         12956 => x"0c",
         12957 => x"04",
         12958 => x"67",
         12959 => x"96",
         12960 => x"52",
         12961 => x"ff",
         12962 => x"84",
         12963 => x"55",
         12964 => x"08",
         12965 => x"38",
         12966 => x"e4",
         12967 => x"0d",
         12968 => x"66",
         12969 => x"d0",
         12970 => x"95",
         12971 => x"b8",
         12972 => x"84",
         12973 => x"e0",
         12974 => x"cf",
         12975 => x"a0",
         12976 => x"55",
         12977 => x"60",
         12978 => x"86",
         12979 => x"90",
         12980 => x"59",
         12981 => x"17",
         12982 => x"2a",
         12983 => x"17",
         12984 => x"2a",
         12985 => x"17",
         12986 => x"2a",
         12987 => x"17",
         12988 => x"81",
         12989 => x"34",
         12990 => x"e1",
         12991 => x"b8",
         12992 => x"b8",
         12993 => x"3d",
         12994 => x"3d",
         12995 => x"5d",
         12996 => x"9a",
         12997 => x"52",
         12998 => x"ff",
         12999 => x"84",
         13000 => x"84",
         13001 => x"30",
         13002 => x"e4",
         13003 => x"25",
         13004 => x"7a",
         13005 => x"38",
         13006 => x"06",
         13007 => x"81",
         13008 => x"30",
         13009 => x"80",
         13010 => x"7b",
         13011 => x"8c",
         13012 => x"76",
         13013 => x"78",
         13014 => x"80",
         13015 => x"11",
         13016 => x"80",
         13017 => x"08",
         13018 => x"f6",
         13019 => x"33",
         13020 => x"74",
         13021 => x"81",
         13022 => x"38",
         13023 => x"53",
         13024 => x"81",
         13025 => x"fe",
         13026 => x"84",
         13027 => x"80",
         13028 => x"ff",
         13029 => x"76",
         13030 => x"78",
         13031 => x"38",
         13032 => x"56",
         13033 => x"56",
         13034 => x"8b",
         13035 => x"56",
         13036 => x"83",
         13037 => x"75",
         13038 => x"83",
         13039 => x"12",
         13040 => x"2b",
         13041 => x"07",
         13042 => x"70",
         13043 => x"2b",
         13044 => x"07",
         13045 => x"5d",
         13046 => x"56",
         13047 => x"e4",
         13048 => x"0d",
         13049 => x"80",
         13050 => x"8e",
         13051 => x"55",
         13052 => x"3f",
         13053 => x"08",
         13054 => x"e4",
         13055 => x"81",
         13056 => x"84",
         13057 => x"06",
         13058 => x"80",
         13059 => x"57",
         13060 => x"77",
         13061 => x"08",
         13062 => x"70",
         13063 => x"33",
         13064 => x"dc",
         13065 => x"59",
         13066 => x"08",
         13067 => x"81",
         13068 => x"38",
         13069 => x"08",
         13070 => x"b4",
         13071 => x"17",
         13072 => x"b8",
         13073 => x"55",
         13074 => x"08",
         13075 => x"38",
         13076 => x"55",
         13077 => x"09",
         13078 => x"a0",
         13079 => x"b4",
         13080 => x"17",
         13081 => x"7a",
         13082 => x"33",
         13083 => x"e2",
         13084 => x"81",
         13085 => x"b8",
         13086 => x"16",
         13087 => x"da",
         13088 => x"b8",
         13089 => x"2e",
         13090 => x"fe",
         13091 => x"52",
         13092 => x"f8",
         13093 => x"b8",
         13094 => x"84",
         13095 => x"fe",
         13096 => x"b8",
         13097 => x"b8",
         13098 => x"5c",
         13099 => x"18",
         13100 => x"1b",
         13101 => x"75",
         13102 => x"81",
         13103 => x"78",
         13104 => x"8b",
         13105 => x"58",
         13106 => x"77",
         13107 => x"f2",
         13108 => x"7b",
         13109 => x"5c",
         13110 => x"a0",
         13111 => x"fc",
         13112 => x"57",
         13113 => x"e1",
         13114 => x"53",
         13115 => x"b4",
         13116 => x"3d",
         13117 => x"eb",
         13118 => x"e4",
         13119 => x"b8",
         13120 => x"a6",
         13121 => x"5d",
         13122 => x"55",
         13123 => x"81",
         13124 => x"ff",
         13125 => x"f4",
         13126 => x"3d",
         13127 => x"70",
         13128 => x"5b",
         13129 => x"9f",
         13130 => x"b7",
         13131 => x"90",
         13132 => x"75",
         13133 => x"81",
         13134 => x"74",
         13135 => x"75",
         13136 => x"83",
         13137 => x"81",
         13138 => x"51",
         13139 => x"83",
         13140 => x"b8",
         13141 => x"9f",
         13142 => x"b8",
         13143 => x"ff",
         13144 => x"76",
         13145 => x"e0",
         13146 => x"f4",
         13147 => x"f4",
         13148 => x"ff",
         13149 => x"58",
         13150 => x"81",
         13151 => x"56",
         13152 => x"99",
         13153 => x"70",
         13154 => x"ff",
         13155 => x"58",
         13156 => x"89",
         13157 => x"2e",
         13158 => x"e9",
         13159 => x"ff",
         13160 => x"81",
         13161 => x"ff",
         13162 => x"f8",
         13163 => x"26",
         13164 => x"81",
         13165 => x"8f",
         13166 => x"2a",
         13167 => x"70",
         13168 => x"34",
         13169 => x"76",
         13170 => x"05",
         13171 => x"1a",
         13172 => x"70",
         13173 => x"ff",
         13174 => x"58",
         13175 => x"26",
         13176 => x"8f",
         13177 => x"86",
         13178 => x"e5",
         13179 => x"79",
         13180 => x"38",
         13181 => x"56",
         13182 => x"33",
         13183 => x"a0",
         13184 => x"06",
         13185 => x"1a",
         13186 => x"38",
         13187 => x"47",
         13188 => x"3d",
         13189 => x"fe",
         13190 => x"84",
         13191 => x"55",
         13192 => x"08",
         13193 => x"38",
         13194 => x"84",
         13195 => x"a1",
         13196 => x"83",
         13197 => x"51",
         13198 => x"84",
         13199 => x"83",
         13200 => x"55",
         13201 => x"38",
         13202 => x"84",
         13203 => x"a1",
         13204 => x"83",
         13205 => x"56",
         13206 => x"81",
         13207 => x"fe",
         13208 => x"84",
         13209 => x"55",
         13210 => x"08",
         13211 => x"79",
         13212 => x"c4",
         13213 => x"7e",
         13214 => x"76",
         13215 => x"58",
         13216 => x"81",
         13217 => x"ff",
         13218 => x"ef",
         13219 => x"81",
         13220 => x"34",
         13221 => x"d9",
         13222 => x"b8",
         13223 => x"74",
         13224 => x"39",
         13225 => x"fe",
         13226 => x"56",
         13227 => x"84",
         13228 => x"84",
         13229 => x"06",
         13230 => x"80",
         13231 => x"2e",
         13232 => x"75",
         13233 => x"76",
         13234 => x"ee",
         13235 => x"b8",
         13236 => x"84",
         13237 => x"75",
         13238 => x"06",
         13239 => x"84",
         13240 => x"b8",
         13241 => x"98",
         13242 => x"80",
         13243 => x"08",
         13244 => x"38",
         13245 => x"55",
         13246 => x"09",
         13247 => x"d7",
         13248 => x"76",
         13249 => x"52",
         13250 => x"51",
         13251 => x"3f",
         13252 => x"08",
         13253 => x"38",
         13254 => x"59",
         13255 => x"0c",
         13256 => x"be",
         13257 => x"17",
         13258 => x"57",
         13259 => x"81",
         13260 => x"9e",
         13261 => x"70",
         13262 => x"07",
         13263 => x"80",
         13264 => x"38",
         13265 => x"79",
         13266 => x"38",
         13267 => x"51",
         13268 => x"3f",
         13269 => x"08",
         13270 => x"e4",
         13271 => x"ff",
         13272 => x"55",
         13273 => x"fd",
         13274 => x"55",
         13275 => x"38",
         13276 => x"55",
         13277 => x"81",
         13278 => x"ff",
         13279 => x"f4",
         13280 => x"88",
         13281 => x"34",
         13282 => x"59",
         13283 => x"70",
         13284 => x"33",
         13285 => x"05",
         13286 => x"15",
         13287 => x"2e",
         13288 => x"76",
         13289 => x"58",
         13290 => x"81",
         13291 => x"ff",
         13292 => x"da",
         13293 => x"39",
         13294 => x"7a",
         13295 => x"81",
         13296 => x"34",
         13297 => x"d7",
         13298 => x"b8",
         13299 => x"fd",
         13300 => x"57",
         13301 => x"81",
         13302 => x"08",
         13303 => x"81",
         13304 => x"fe",
         13305 => x"84",
         13306 => x"79",
         13307 => x"06",
         13308 => x"84",
         13309 => x"83",
         13310 => x"18",
         13311 => x"08",
         13312 => x"a0",
         13313 => x"8a",
         13314 => x"33",
         13315 => x"2e",
         13316 => x"b8",
         13317 => x"fd",
         13318 => x"5a",
         13319 => x"51",
         13320 => x"3f",
         13321 => x"08",
         13322 => x"e4",
         13323 => x"fd",
         13324 => x"ae",
         13325 => x"58",
         13326 => x"2e",
         13327 => x"fe",
         13328 => x"54",
         13329 => x"a0",
         13330 => x"53",
         13331 => x"18",
         13332 => x"d3",
         13333 => x"a9",
         13334 => x"0d",
         13335 => x"88",
         13336 => x"05",
         13337 => x"57",
         13338 => x"80",
         13339 => x"76",
         13340 => x"80",
         13341 => x"74",
         13342 => x"80",
         13343 => x"86",
         13344 => x"18",
         13345 => x"78",
         13346 => x"c2",
         13347 => x"73",
         13348 => x"a5",
         13349 => x"33",
         13350 => x"9d",
         13351 => x"2e",
         13352 => x"8c",
         13353 => x"9c",
         13354 => x"33",
         13355 => x"81",
         13356 => x"74",
         13357 => x"8c",
         13358 => x"11",
         13359 => x"2b",
         13360 => x"54",
         13361 => x"fd",
         13362 => x"ff",
         13363 => x"70",
         13364 => x"07",
         13365 => x"b8",
         13366 => x"90",
         13367 => x"42",
         13368 => x"58",
         13369 => x"88",
         13370 => x"08",
         13371 => x"38",
         13372 => x"78",
         13373 => x"59",
         13374 => x"51",
         13375 => x"3f",
         13376 => x"55",
         13377 => x"08",
         13378 => x"38",
         13379 => x"b8",
         13380 => x"2e",
         13381 => x"84",
         13382 => x"ff",
         13383 => x"38",
         13384 => x"08",
         13385 => x"81",
         13386 => x"7d",
         13387 => x"74",
         13388 => x"81",
         13389 => x"87",
         13390 => x"73",
         13391 => x"0c",
         13392 => x"04",
         13393 => x"b8",
         13394 => x"3d",
         13395 => x"15",
         13396 => x"d0",
         13397 => x"b8",
         13398 => x"06",
         13399 => x"ad",
         13400 => x"08",
         13401 => x"a7",
         13402 => x"2e",
         13403 => x"7a",
         13404 => x"7c",
         13405 => x"38",
         13406 => x"74",
         13407 => x"e6",
         13408 => x"77",
         13409 => x"fe",
         13410 => x"84",
         13411 => x"56",
         13412 => x"08",
         13413 => x"77",
         13414 => x"17",
         13415 => x"74",
         13416 => x"7e",
         13417 => x"55",
         13418 => x"ff",
         13419 => x"88",
         13420 => x"8c",
         13421 => x"17",
         13422 => x"07",
         13423 => x"18",
         13424 => x"08",
         13425 => x"16",
         13426 => x"76",
         13427 => x"e9",
         13428 => x"31",
         13429 => x"84",
         13430 => x"07",
         13431 => x"16",
         13432 => x"fe",
         13433 => x"54",
         13434 => x"74",
         13435 => x"fe",
         13436 => x"54",
         13437 => x"81",
         13438 => x"39",
         13439 => x"ff",
         13440 => x"b8",
         13441 => x"3d",
         13442 => x"08",
         13443 => x"02",
         13444 => x"87",
         13445 => x"42",
         13446 => x"a2",
         13447 => x"5f",
         13448 => x"80",
         13449 => x"38",
         13450 => x"05",
         13451 => x"9f",
         13452 => x"75",
         13453 => x"9b",
         13454 => x"38",
         13455 => x"85",
         13456 => x"d0",
         13457 => x"80",
         13458 => x"e5",
         13459 => x"10",
         13460 => x"05",
         13461 => x"5a",
         13462 => x"84",
         13463 => x"34",
         13464 => x"b8",
         13465 => x"84",
         13466 => x"33",
         13467 => x"81",
         13468 => x"fe",
         13469 => x"84",
         13470 => x"81",
         13471 => x"81",
         13472 => x"83",
         13473 => x"ab",
         13474 => x"2a",
         13475 => x"8a",
         13476 => x"9f",
         13477 => x"fc",
         13478 => x"52",
         13479 => x"d0",
         13480 => x"b8",
         13481 => x"98",
         13482 => x"74",
         13483 => x"90",
         13484 => x"80",
         13485 => x"88",
         13486 => x"75",
         13487 => x"83",
         13488 => x"80",
         13489 => x"84",
         13490 => x"83",
         13491 => x"81",
         13492 => x"83",
         13493 => x"1f",
         13494 => x"74",
         13495 => x"7e",
         13496 => x"3d",
         13497 => x"70",
         13498 => x"59",
         13499 => x"60",
         13500 => x"ab",
         13501 => x"70",
         13502 => x"07",
         13503 => x"57",
         13504 => x"38",
         13505 => x"84",
         13506 => x"54",
         13507 => x"52",
         13508 => x"cd",
         13509 => x"57",
         13510 => x"08",
         13511 => x"60",
         13512 => x"33",
         13513 => x"05",
         13514 => x"2b",
         13515 => x"8e",
         13516 => x"d4",
         13517 => x"81",
         13518 => x"38",
         13519 => x"61",
         13520 => x"11",
         13521 => x"62",
         13522 => x"e7",
         13523 => x"18",
         13524 => x"82",
         13525 => x"90",
         13526 => x"2b",
         13527 => x"33",
         13528 => x"88",
         13529 => x"71",
         13530 => x"1f",
         13531 => x"82",
         13532 => x"90",
         13533 => x"2b",
         13534 => x"33",
         13535 => x"88",
         13536 => x"71",
         13537 => x"3d",
         13538 => x"3d",
         13539 => x"0c",
         13540 => x"45",
         13541 => x"5a",
         13542 => x"8e",
         13543 => x"79",
         13544 => x"38",
         13545 => x"81",
         13546 => x"87",
         13547 => x"2a",
         13548 => x"45",
         13549 => x"2e",
         13550 => x"61",
         13551 => x"64",
         13552 => x"38",
         13553 => x"47",
         13554 => x"38",
         13555 => x"30",
         13556 => x"7a",
         13557 => x"2e",
         13558 => x"7a",
         13559 => x"8c",
         13560 => x"0b",
         13561 => x"22",
         13562 => x"80",
         13563 => x"74",
         13564 => x"38",
         13565 => x"56",
         13566 => x"17",
         13567 => x"57",
         13568 => x"2e",
         13569 => x"75",
         13570 => x"77",
         13571 => x"fd",
         13572 => x"84",
         13573 => x"10",
         13574 => x"84",
         13575 => x"9f",
         13576 => x"38",
         13577 => x"b8",
         13578 => x"84",
         13579 => x"05",
         13580 => x"2a",
         13581 => x"4c",
         13582 => x"15",
         13583 => x"81",
         13584 => x"7b",
         13585 => x"68",
         13586 => x"ff",
         13587 => x"06",
         13588 => x"4e",
         13589 => x"83",
         13590 => x"38",
         13591 => x"77",
         13592 => x"70",
         13593 => x"57",
         13594 => x"82",
         13595 => x"7c",
         13596 => x"78",
         13597 => x"31",
         13598 => x"80",
         13599 => x"b8",
         13600 => x"62",
         13601 => x"f6",
         13602 => x"2e",
         13603 => x"82",
         13604 => x"ff",
         13605 => x"b8",
         13606 => x"82",
         13607 => x"89",
         13608 => x"18",
         13609 => x"c0",
         13610 => x"38",
         13611 => x"a3",
         13612 => x"76",
         13613 => x"0c",
         13614 => x"84",
         13615 => x"04",
         13616 => x"fe",
         13617 => x"84",
         13618 => x"9f",
         13619 => x"b8",
         13620 => x"7c",
         13621 => x"70",
         13622 => x"57",
         13623 => x"89",
         13624 => x"82",
         13625 => x"ff",
         13626 => x"5d",
         13627 => x"2e",
         13628 => x"80",
         13629 => x"d4",
         13630 => x"08",
         13631 => x"7a",
         13632 => x"5c",
         13633 => x"81",
         13634 => x"ff",
         13635 => x"59",
         13636 => x"26",
         13637 => x"17",
         13638 => x"06",
         13639 => x"9f",
         13640 => x"99",
         13641 => x"e0",
         13642 => x"ff",
         13643 => x"76",
         13644 => x"2a",
         13645 => x"78",
         13646 => x"06",
         13647 => x"ff",
         13648 => x"7a",
         13649 => x"70",
         13650 => x"2a",
         13651 => x"4a",
         13652 => x"2e",
         13653 => x"81",
         13654 => x"5f",
         13655 => x"25",
         13656 => x"7f",
         13657 => x"39",
         13658 => x"05",
         13659 => x"79",
         13660 => x"dd",
         13661 => x"84",
         13662 => x"fe",
         13663 => x"83",
         13664 => x"84",
         13665 => x"40",
         13666 => x"38",
         13667 => x"55",
         13668 => x"75",
         13669 => x"38",
         13670 => x"59",
         13671 => x"81",
         13672 => x"39",
         13673 => x"ff",
         13674 => x"7a",
         13675 => x"56",
         13676 => x"61",
         13677 => x"93",
         13678 => x"2e",
         13679 => x"82",
         13680 => x"4a",
         13681 => x"8b",
         13682 => x"e4",
         13683 => x"26",
         13684 => x"8b",
         13685 => x"5b",
         13686 => x"27",
         13687 => x"8e",
         13688 => x"b8",
         13689 => x"3d",
         13690 => x"f0",
         13691 => x"55",
         13692 => x"86",
         13693 => x"f5",
         13694 => x"38",
         13695 => x"5b",
         13696 => x"fd",
         13697 => x"80",
         13698 => x"80",
         13699 => x"05",
         13700 => x"15",
         13701 => x"38",
         13702 => x"e4",
         13703 => x"55",
         13704 => x"05",
         13705 => x"70",
         13706 => x"34",
         13707 => x"74",
         13708 => x"8b",
         13709 => x"65",
         13710 => x"8c",
         13711 => x"61",
         13712 => x"7b",
         13713 => x"06",
         13714 => x"8e",
         13715 => x"88",
         13716 => x"61",
         13717 => x"81",
         13718 => x"34",
         13719 => x"70",
         13720 => x"80",
         13721 => x"34",
         13722 => x"82",
         13723 => x"61",
         13724 => x"6c",
         13725 => x"ff",
         13726 => x"ad",
         13727 => x"ff",
         13728 => x"74",
         13729 => x"34",
         13730 => x"4c",
         13731 => x"05",
         13732 => x"95",
         13733 => x"61",
         13734 => x"80",
         13735 => x"34",
         13736 => x"05",
         13737 => x"9b",
         13738 => x"61",
         13739 => x"7e",
         13740 => x"67",
         13741 => x"34",
         13742 => x"4c",
         13743 => x"05",
         13744 => x"2a",
         13745 => x"0c",
         13746 => x"08",
         13747 => x"34",
         13748 => x"85",
         13749 => x"61",
         13750 => x"80",
         13751 => x"34",
         13752 => x"05",
         13753 => x"61",
         13754 => x"7c",
         13755 => x"06",
         13756 => x"96",
         13757 => x"88",
         13758 => x"61",
         13759 => x"ff",
         13760 => x"05",
         13761 => x"a6",
         13762 => x"61",
         13763 => x"e4",
         13764 => x"55",
         13765 => x"05",
         13766 => x"70",
         13767 => x"34",
         13768 => x"74",
         13769 => x"83",
         13770 => x"80",
         13771 => x"60",
         13772 => x"4b",
         13773 => x"34",
         13774 => x"53",
         13775 => x"51",
         13776 => x"3f",
         13777 => x"b8",
         13778 => x"e7",
         13779 => x"5c",
         13780 => x"87",
         13781 => x"61",
         13782 => x"76",
         13783 => x"58",
         13784 => x"55",
         13785 => x"63",
         13786 => x"62",
         13787 => x"c0",
         13788 => x"ff",
         13789 => x"81",
         13790 => x"f8",
         13791 => x"34",
         13792 => x"7c",
         13793 => x"64",
         13794 => x"46",
         13795 => x"2a",
         13796 => x"70",
         13797 => x"34",
         13798 => x"56",
         13799 => x"7c",
         13800 => x"76",
         13801 => x"38",
         13802 => x"54",
         13803 => x"52",
         13804 => x"c5",
         13805 => x"b8",
         13806 => x"e6",
         13807 => x"61",
         13808 => x"76",
         13809 => x"58",
         13810 => x"55",
         13811 => x"78",
         13812 => x"31",
         13813 => x"c9",
         13814 => x"05",
         13815 => x"2e",
         13816 => x"77",
         13817 => x"2e",
         13818 => x"56",
         13819 => x"66",
         13820 => x"75",
         13821 => x"7a",
         13822 => x"79",
         13823 => x"d2",
         13824 => x"e4",
         13825 => x"38",
         13826 => x"76",
         13827 => x"75",
         13828 => x"58",
         13829 => x"93",
         13830 => x"6c",
         13831 => x"26",
         13832 => x"58",
         13833 => x"83",
         13834 => x"7d",
         13835 => x"61",
         13836 => x"06",
         13837 => x"b3",
         13838 => x"61",
         13839 => x"75",
         13840 => x"57",
         13841 => x"59",
         13842 => x"80",
         13843 => x"ff",
         13844 => x"60",
         13845 => x"47",
         13846 => x"81",
         13847 => x"34",
         13848 => x"05",
         13849 => x"83",
         13850 => x"67",
         13851 => x"6c",
         13852 => x"c1",
         13853 => x"51",
         13854 => x"3f",
         13855 => x"05",
         13856 => x"e4",
         13857 => x"bf",
         13858 => x"67",
         13859 => x"84",
         13860 => x"67",
         13861 => x"7e",
         13862 => x"05",
         13863 => x"83",
         13864 => x"6b",
         13865 => x"05",
         13866 => x"f0",
         13867 => x"c9",
         13868 => x"61",
         13869 => x"34",
         13870 => x"45",
         13871 => x"cb",
         13872 => x"90",
         13873 => x"61",
         13874 => x"34",
         13875 => x"5f",
         13876 => x"cd",
         13877 => x"54",
         13878 => x"52",
         13879 => x"c2",
         13880 => x"57",
         13881 => x"08",
         13882 => x"80",
         13883 => x"79",
         13884 => x"dd",
         13885 => x"84",
         13886 => x"f7",
         13887 => x"b8",
         13888 => x"b8",
         13889 => x"3d",
         13890 => x"f0",
         13891 => x"55",
         13892 => x"74",
         13893 => x"45",
         13894 => x"39",
         13895 => x"78",
         13896 => x"81",
         13897 => x"98",
         13898 => x"74",
         13899 => x"38",
         13900 => x"98",
         13901 => x"98",
         13902 => x"82",
         13903 => x"57",
         13904 => x"80",
         13905 => x"76",
         13906 => x"38",
         13907 => x"51",
         13908 => x"3f",
         13909 => x"08",
         13910 => x"87",
         13911 => x"2a",
         13912 => x"5c",
         13913 => x"b8",
         13914 => x"80",
         13915 => x"47",
         13916 => x"0a",
         13917 => x"cb",
         13918 => x"f8",
         13919 => x"b8",
         13920 => x"ff",
         13921 => x"e6",
         13922 => x"d3",
         13923 => x"2a",
         13924 => x"bf",
         13925 => x"f8",
         13926 => x"81",
         13927 => x"80",
         13928 => x"38",
         13929 => x"ab",
         13930 => x"a0",
         13931 => x"88",
         13932 => x"61",
         13933 => x"75",
         13934 => x"7a",
         13935 => x"34",
         13936 => x"57",
         13937 => x"05",
         13938 => x"39",
         13939 => x"c3",
         13940 => x"61",
         13941 => x"34",
         13942 => x"c5",
         13943 => x"cc",
         13944 => x"05",
         13945 => x"a4",
         13946 => x"88",
         13947 => x"61",
         13948 => x"7c",
         13949 => x"78",
         13950 => x"34",
         13951 => x"56",
         13952 => x"05",
         13953 => x"ac",
         13954 => x"61",
         13955 => x"80",
         13956 => x"34",
         13957 => x"05",
         13958 => x"b0",
         13959 => x"61",
         13960 => x"86",
         13961 => x"34",
         13962 => x"05",
         13963 => x"61",
         13964 => x"34",
         13965 => x"c2",
         13966 => x"61",
         13967 => x"83",
         13968 => x"57",
         13969 => x"81",
         13970 => x"76",
         13971 => x"58",
         13972 => x"55",
         13973 => x"f9",
         13974 => x"70",
         13975 => x"33",
         13976 => x"05",
         13977 => x"15",
         13978 => x"38",
         13979 => x"81",
         13980 => x"60",
         13981 => x"fe",
         13982 => x"81",
         13983 => x"e4",
         13984 => x"38",
         13985 => x"61",
         13986 => x"62",
         13987 => x"34",
         13988 => x"b8",
         13989 => x"60",
         13990 => x"fe",
         13991 => x"fc",
         13992 => x"0b",
         13993 => x"0c",
         13994 => x"84",
         13995 => x"04",
         13996 => x"7b",
         13997 => x"70",
         13998 => x"34",
         13999 => x"81",
         14000 => x"ff",
         14001 => x"61",
         14002 => x"ff",
         14003 => x"34",
         14004 => x"05",
         14005 => x"87",
         14006 => x"61",
         14007 => x"ff",
         14008 => x"34",
         14009 => x"05",
         14010 => x"34",
         14011 => x"b1",
         14012 => x"86",
         14013 => x"52",
         14014 => x"be",
         14015 => x"80",
         14016 => x"80",
         14017 => x"05",
         14018 => x"17",
         14019 => x"38",
         14020 => x"d2",
         14021 => x"05",
         14022 => x"55",
         14023 => x"70",
         14024 => x"34",
         14025 => x"70",
         14026 => x"34",
         14027 => x"34",
         14028 => x"83",
         14029 => x"80",
         14030 => x"e5",
         14031 => x"c1",
         14032 => x"05",
         14033 => x"61",
         14034 => x"34",
         14035 => x"5b",
         14036 => x"e8",
         14037 => x"88",
         14038 => x"61",
         14039 => x"34",
         14040 => x"56",
         14041 => x"ea",
         14042 => x"98",
         14043 => x"61",
         14044 => x"34",
         14045 => x"ec",
         14046 => x"61",
         14047 => x"34",
         14048 => x"ee",
         14049 => x"61",
         14050 => x"34",
         14051 => x"34",
         14052 => x"34",
         14053 => x"1f",
         14054 => x"79",
         14055 => x"b2",
         14056 => x"81",
         14057 => x"52",
         14058 => x"bd",
         14059 => x"61",
         14060 => x"a6",
         14061 => x"0d",
         14062 => x"5b",
         14063 => x"ff",
         14064 => x"57",
         14065 => x"b8",
         14066 => x"59",
         14067 => x"05",
         14068 => x"78",
         14069 => x"ff",
         14070 => x"7b",
         14071 => x"81",
         14072 => x"8d",
         14073 => x"74",
         14074 => x"38",
         14075 => x"81",
         14076 => x"81",
         14077 => x"8a",
         14078 => x"77",
         14079 => x"38",
         14080 => x"7a",
         14081 => x"38",
         14082 => x"84",
         14083 => x"8e",
         14084 => x"f7",
         14085 => x"02",
         14086 => x"05",
         14087 => x"77",
         14088 => x"d5",
         14089 => x"08",
         14090 => x"24",
         14091 => x"17",
         14092 => x"8c",
         14093 => x"77",
         14094 => x"16",
         14095 => x"24",
         14096 => x"84",
         14097 => x"19",
         14098 => x"8b",
         14099 => x"8b",
         14100 => x"54",
         14101 => x"17",
         14102 => x"51",
         14103 => x"3f",
         14104 => x"70",
         14105 => x"07",
         14106 => x"30",
         14107 => x"81",
         14108 => x"0c",
         14109 => x"d3",
         14110 => x"76",
         14111 => x"3f",
         14112 => x"e3",
         14113 => x"80",
         14114 => x"8d",
         14115 => x"80",
         14116 => x"55",
         14117 => x"81",
         14118 => x"ff",
         14119 => x"f4",
         14120 => x"08",
         14121 => x"8a",
         14122 => x"38",
         14123 => x"76",
         14124 => x"38",
         14125 => x"8c",
         14126 => x"77",
         14127 => x"16",
         14128 => x"24",
         14129 => x"84",
         14130 => x"19",
         14131 => x"7c",
         14132 => x"24",
         14133 => x"3d",
         14134 => x"55",
         14135 => x"05",
         14136 => x"51",
         14137 => x"3f",
         14138 => x"08",
         14139 => x"7a",
         14140 => x"ff",
         14141 => x"e4",
         14142 => x"0d",
         14143 => x"ff",
         14144 => x"75",
         14145 => x"52",
         14146 => x"ff",
         14147 => x"74",
         14148 => x"30",
         14149 => x"9f",
         14150 => x"52",
         14151 => x"ff",
         14152 => x"52",
         14153 => x"eb",
         14154 => x"39",
         14155 => x"e4",
         14156 => x"0d",
         14157 => x"0d",
         14158 => x"05",
         14159 => x"52",
         14160 => x"72",
         14161 => x"90",
         14162 => x"ff",
         14163 => x"71",
         14164 => x"0c",
         14165 => x"04",
         14166 => x"73",
         14167 => x"83",
         14168 => x"81",
         14169 => x"73",
         14170 => x"38",
         14171 => x"22",
         14172 => x"2e",
         14173 => x"12",
         14174 => x"ff",
         14175 => x"71",
         14176 => x"8d",
         14177 => x"83",
         14178 => x"70",
         14179 => x"e1",
         14180 => x"12",
         14181 => x"06",
         14182 => x"0c",
         14183 => x"0d",
         14184 => x"0d",
         14185 => x"22",
         14186 => x"96",
         14187 => x"51",
         14188 => x"80",
         14189 => x"38",
         14190 => x"84",
         14191 => x"84",
         14192 => x"71",
         14193 => x"09",
         14194 => x"38",
         14195 => x"26",
         14196 => x"10",
         14197 => x"05",
         14198 => x"b8",
         14199 => x"84",
         14200 => x"fb",
         14201 => x"51",
         14202 => x"ff",
         14203 => x"38",
         14204 => x"ff",
         14205 => x"a8",
         14206 => x"9f",
         14207 => x"d9",
         14208 => x"82",
         14209 => x"75",
         14210 => x"80",
         14211 => x"26",
         14212 => x"53",
         14213 => x"38",
         14214 => x"05",
         14215 => x"71",
         14216 => x"56",
         14217 => x"70",
         14218 => x"70",
         14219 => x"38",
         14220 => x"73",
         14221 => x"70",
         14222 => x"22",
         14223 => x"70",
         14224 => x"79",
         14225 => x"55",
         14226 => x"2e",
         14227 => x"51",
         14228 => x"e4",
         14229 => x"0d",
         14230 => x"9c",
         14231 => x"39",
         14232 => x"ea",
         14233 => x"10",
         14234 => x"05",
         14235 => x"04",
         14236 => x"70",
         14237 => x"06",
         14238 => x"51",
         14239 => x"b0",
         14240 => x"ff",
         14241 => x"51",
         14242 => x"16",
         14243 => x"ff",
         14244 => x"e6",
         14245 => x"70",
         14246 => x"06",
         14247 => x"39",
         14248 => x"83",
         14249 => x"57",
         14250 => x"e0",
         14251 => x"ff",
         14252 => x"51",
         14253 => x"16",
         14254 => x"ff",
         14255 => x"ff",
         14256 => x"73",
         14257 => x"76",
         14258 => x"83",
         14259 => x"58",
         14260 => x"a6",
         14261 => x"31",
         14262 => x"70",
         14263 => x"fe",
         14264 => x"00",
         14265 => x"ff",
         14266 => x"ff",
         14267 => x"00",
         14268 => x"ff",
         14269 => x"19",
         14270 => x"19",
         14271 => x"19",
         14272 => x"19",
         14273 => x"19",
         14274 => x"19",
         14275 => x"19",
         14276 => x"19",
         14277 => x"19",
         14278 => x"19",
         14279 => x"19",
         14280 => x"19",
         14281 => x"19",
         14282 => x"18",
         14283 => x"18",
         14284 => x"18",
         14285 => x"18",
         14286 => x"18",
         14287 => x"18",
         14288 => x"18",
         14289 => x"1e",
         14290 => x"1f",
         14291 => x"1f",
         14292 => x"1f",
         14293 => x"1f",
         14294 => x"1f",
         14295 => x"1f",
         14296 => x"1f",
         14297 => x"1f",
         14298 => x"1f",
         14299 => x"1f",
         14300 => x"1f",
         14301 => x"1f",
         14302 => x"1f",
         14303 => x"1f",
         14304 => x"1f",
         14305 => x"1f",
         14306 => x"1f",
         14307 => x"1f",
         14308 => x"1f",
         14309 => x"1f",
         14310 => x"1f",
         14311 => x"1f",
         14312 => x"1f",
         14313 => x"1f",
         14314 => x"1f",
         14315 => x"1f",
         14316 => x"1f",
         14317 => x"1f",
         14318 => x"1f",
         14319 => x"1f",
         14320 => x"1f",
         14321 => x"1f",
         14322 => x"1f",
         14323 => x"1f",
         14324 => x"1f",
         14325 => x"1f",
         14326 => x"1f",
         14327 => x"1f",
         14328 => x"1f",
         14329 => x"1f",
         14330 => x"1f",
         14331 => x"1f",
         14332 => x"24",
         14333 => x"1f",
         14334 => x"1f",
         14335 => x"1f",
         14336 => x"1f",
         14337 => x"1f",
         14338 => x"1f",
         14339 => x"1f",
         14340 => x"1f",
         14341 => x"1f",
         14342 => x"1f",
         14343 => x"1f",
         14344 => x"1f",
         14345 => x"1f",
         14346 => x"1f",
         14347 => x"1f",
         14348 => x"1f",
         14349 => x"24",
         14350 => x"23",
         14351 => x"1f",
         14352 => x"22",
         14353 => x"24",
         14354 => x"23",
         14355 => x"22",
         14356 => x"21",
         14357 => x"1f",
         14358 => x"1f",
         14359 => x"1f",
         14360 => x"1f",
         14361 => x"1f",
         14362 => x"1f",
         14363 => x"1f",
         14364 => x"1f",
         14365 => x"1f",
         14366 => x"1f",
         14367 => x"1f",
         14368 => x"1f",
         14369 => x"1f",
         14370 => x"1f",
         14371 => x"1f",
         14372 => x"1f",
         14373 => x"1f",
         14374 => x"1f",
         14375 => x"1f",
         14376 => x"1f",
         14377 => x"1f",
         14378 => x"1f",
         14379 => x"1f",
         14380 => x"1f",
         14381 => x"1f",
         14382 => x"1f",
         14383 => x"1f",
         14384 => x"1f",
         14385 => x"1f",
         14386 => x"1f",
         14387 => x"1f",
         14388 => x"1f",
         14389 => x"1f",
         14390 => x"1f",
         14391 => x"1f",
         14392 => x"1f",
         14393 => x"1f",
         14394 => x"1f",
         14395 => x"1f",
         14396 => x"1f",
         14397 => x"1f",
         14398 => x"1f",
         14399 => x"1f",
         14400 => x"1f",
         14401 => x"1f",
         14402 => x"1f",
         14403 => x"1f",
         14404 => x"1f",
         14405 => x"1f",
         14406 => x"1f",
         14407 => x"1f",
         14408 => x"1f",
         14409 => x"21",
         14410 => x"21",
         14411 => x"1f",
         14412 => x"1f",
         14413 => x"1f",
         14414 => x"1f",
         14415 => x"1f",
         14416 => x"1f",
         14417 => x"1f",
         14418 => x"1f",
         14419 => x"21",
         14420 => x"21",
         14421 => x"1f",
         14422 => x"21",
         14423 => x"1f",
         14424 => x"21",
         14425 => x"21",
         14426 => x"21",
         14427 => x"32",
         14428 => x"32",
         14429 => x"32",
         14430 => x"32",
         14431 => x"32",
         14432 => x"32",
         14433 => x"3b",
         14434 => x"3a",
         14435 => x"38",
         14436 => x"36",
         14437 => x"3a",
         14438 => x"34",
         14439 => x"37",
         14440 => x"36",
         14441 => x"39",
         14442 => x"36",
         14443 => x"37",
         14444 => x"39",
         14445 => x"34",
         14446 => x"38",
         14447 => x"37",
         14448 => x"37",
         14449 => x"34",
         14450 => x"34",
         14451 => x"37",
         14452 => x"36",
         14453 => x"36",
         14454 => x"36",
         14455 => x"46",
         14456 => x"46",
         14457 => x"46",
         14458 => x"46",
         14459 => x"46",
         14460 => x"46",
         14461 => x"46",
         14462 => x"47",
         14463 => x"47",
         14464 => x"47",
         14465 => x"47",
         14466 => x"47",
         14467 => x"47",
         14468 => x"47",
         14469 => x"47",
         14470 => x"47",
         14471 => x"47",
         14472 => x"47",
         14473 => x"47",
         14474 => x"47",
         14475 => x"47",
         14476 => x"47",
         14477 => x"47",
         14478 => x"47",
         14479 => x"47",
         14480 => x"47",
         14481 => x"47",
         14482 => x"47",
         14483 => x"47",
         14484 => x"47",
         14485 => x"47",
         14486 => x"47",
         14487 => x"47",
         14488 => x"47",
         14489 => x"47",
         14490 => x"47",
         14491 => x"47",
         14492 => x"48",
         14493 => x"48",
         14494 => x"48",
         14495 => x"48",
         14496 => x"47",
         14497 => x"48",
         14498 => x"48",
         14499 => x"47",
         14500 => x"47",
         14501 => x"47",
         14502 => x"47",
         14503 => x"48",
         14504 => x"47",
         14505 => x"47",
         14506 => x"47",
         14507 => x"47",
         14508 => x"47",
         14509 => x"47",
         14510 => x"47",
         14511 => x"47",
         14512 => x"53",
         14513 => x"55",
         14514 => x"55",
         14515 => x"54",
         14516 => x"54",
         14517 => x"54",
         14518 => x"54",
         14519 => x"55",
         14520 => x"52",
         14521 => x"55",
         14522 => x"57",
         14523 => x"52",
         14524 => x"52",
         14525 => x"52",
         14526 => x"52",
         14527 => x"52",
         14528 => x"52",
         14529 => x"55",
         14530 => x"57",
         14531 => x"56",
         14532 => x"52",
         14533 => x"52",
         14534 => x"52",
         14535 => x"52",
         14536 => x"52",
         14537 => x"52",
         14538 => x"52",
         14539 => x"52",
         14540 => x"52",
         14541 => x"52",
         14542 => x"52",
         14543 => x"52",
         14544 => x"52",
         14545 => x"52",
         14546 => x"52",
         14547 => x"52",
         14548 => x"52",
         14549 => x"52",
         14550 => x"52",
         14551 => x"55",
         14552 => x"52",
         14553 => x"52",
         14554 => x"52",
         14555 => x"54",
         14556 => x"53",
         14557 => x"53",
         14558 => x"52",
         14559 => x"52",
         14560 => x"52",
         14561 => x"52",
         14562 => x"53",
         14563 => x"52",
         14564 => x"53",
         14565 => x"59",
         14566 => x"59",
         14567 => x"59",
         14568 => x"59",
         14569 => x"59",
         14570 => x"59",
         14571 => x"59",
         14572 => x"58",
         14573 => x"59",
         14574 => x"59",
         14575 => x"59",
         14576 => x"59",
         14577 => x"59",
         14578 => x"59",
         14579 => x"59",
         14580 => x"59",
         14581 => x"59",
         14582 => x"59",
         14583 => x"59",
         14584 => x"59",
         14585 => x"59",
         14586 => x"59",
         14587 => x"59",
         14588 => x"59",
         14589 => x"59",
         14590 => x"59",
         14591 => x"59",
         14592 => x"59",
         14593 => x"59",
         14594 => x"59",
         14595 => x"59",
         14596 => x"59",
         14597 => x"59",
         14598 => x"59",
         14599 => x"59",
         14600 => x"5a",
         14601 => x"5a",
         14602 => x"5a",
         14603 => x"59",
         14604 => x"5a",
         14605 => x"5a",
         14606 => x"5a",
         14607 => x"5a",
         14608 => x"5a",
         14609 => x"59",
         14610 => x"59",
         14611 => x"59",
         14612 => x"59",
         14613 => x"59",
         14614 => x"59",
         14615 => x"63",
         14616 => x"61",
         14617 => x"61",
         14618 => x"61",
         14619 => x"61",
         14620 => x"61",
         14621 => x"61",
         14622 => x"61",
         14623 => x"61",
         14624 => x"61",
         14625 => x"61",
         14626 => x"61",
         14627 => x"61",
         14628 => x"61",
         14629 => x"5e",
         14630 => x"61",
         14631 => x"61",
         14632 => x"61",
         14633 => x"61",
         14634 => x"61",
         14635 => x"61",
         14636 => x"63",
         14637 => x"61",
         14638 => x"61",
         14639 => x"63",
         14640 => x"61",
         14641 => x"63",
         14642 => x"5e",
         14643 => x"63",
         14644 => x"de",
         14645 => x"de",
         14646 => x"de",
         14647 => x"de",
         14648 => x"de",
         14649 => x"de",
         14650 => x"de",
         14651 => x"de",
         14652 => x"de",
         14653 => x"0e",
         14654 => x"0b",
         14655 => x"0b",
         14656 => x"0f",
         14657 => x"0b",
         14658 => x"0b",
         14659 => x"0b",
         14660 => x"0b",
         14661 => x"0b",
         14662 => x"0b",
         14663 => x"0b",
         14664 => x"0d",
         14665 => x"0b",
         14666 => x"0f",
         14667 => x"0f",
         14668 => x"0b",
         14669 => x"0b",
         14670 => x"0b",
         14671 => x"0b",
         14672 => x"0b",
         14673 => x"0b",
         14674 => x"0b",
         14675 => x"0b",
         14676 => x"0b",
         14677 => x"0b",
         14678 => x"0b",
         14679 => x"0b",
         14680 => x"0b",
         14681 => x"0b",
         14682 => x"0b",
         14683 => x"0b",
         14684 => x"0b",
         14685 => x"0b",
         14686 => x"0b",
         14687 => x"0b",
         14688 => x"0b",
         14689 => x"0b",
         14690 => x"0b",
         14691 => x"0b",
         14692 => x"0b",
         14693 => x"0b",
         14694 => x"0b",
         14695 => x"0b",
         14696 => x"0b",
         14697 => x"0b",
         14698 => x"0b",
         14699 => x"0b",
         14700 => x"0b",
         14701 => x"0b",
         14702 => x"0b",
         14703 => x"0b",
         14704 => x"0f",
         14705 => x"0b",
         14706 => x"0b",
         14707 => x"0b",
         14708 => x"0b",
         14709 => x"0e",
         14710 => x"0b",
         14711 => x"0b",
         14712 => x"0b",
         14713 => x"0b",
         14714 => x"0b",
         14715 => x"0b",
         14716 => x"0b",
         14717 => x"0b",
         14718 => x"0b",
         14719 => x"0b",
         14720 => x"0e",
         14721 => x"0e",
         14722 => x"0e",
         14723 => x"0e",
         14724 => x"0e",
         14725 => x"0b",
         14726 => x"0e",
         14727 => x"0b",
         14728 => x"0b",
         14729 => x"0e",
         14730 => x"0b",
         14731 => x"0b",
         14732 => x"0c",
         14733 => x"0e",
         14734 => x"0b",
         14735 => x"0b",
         14736 => x"0f",
         14737 => x"0b",
         14738 => x"0c",
         14739 => x"0b",
         14740 => x"0b",
         14741 => x"0e",
         14742 => x"6e",
         14743 => x"00",
         14744 => x"6f",
         14745 => x"00",
         14746 => x"6e",
         14747 => x"00",
         14748 => x"6f",
         14749 => x"00",
         14750 => x"78",
         14751 => x"00",
         14752 => x"6c",
         14753 => x"00",
         14754 => x"6f",
         14755 => x"00",
         14756 => x"69",
         14757 => x"00",
         14758 => x"75",
         14759 => x"00",
         14760 => x"62",
         14761 => x"68",
         14762 => x"77",
         14763 => x"64",
         14764 => x"65",
         14765 => x"64",
         14766 => x"65",
         14767 => x"6c",
         14768 => x"00",
         14769 => x"70",
         14770 => x"73",
         14771 => x"74",
         14772 => x"73",
         14773 => x"00",
         14774 => x"66",
         14775 => x"00",
         14776 => x"73",
         14777 => x"00",
         14778 => x"73",
         14779 => x"30",
         14780 => x"61",
         14781 => x"00",
         14782 => x"61",
         14783 => x"00",
         14784 => x"6c",
         14785 => x"00",
         14786 => x"00",
         14787 => x"6b",
         14788 => x"6e",
         14789 => x"72",
         14790 => x"00",
         14791 => x"72",
         14792 => x"74",
         14793 => x"20",
         14794 => x"6f",
         14795 => x"63",
         14796 => x"00",
         14797 => x"6f",
         14798 => x"6e",
         14799 => x"70",
         14800 => x"66",
         14801 => x"73",
         14802 => x"00",
         14803 => x"73",
         14804 => x"69",
         14805 => x"6e",
         14806 => x"65",
         14807 => x"79",
         14808 => x"00",
         14809 => x"6c",
         14810 => x"73",
         14811 => x"63",
         14812 => x"2e",
         14813 => x"6d",
         14814 => x"74",
         14815 => x"70",
         14816 => x"74",
         14817 => x"20",
         14818 => x"63",
         14819 => x"65",
         14820 => x"00",
         14821 => x"72",
         14822 => x"20",
         14823 => x"72",
         14824 => x"2e",
         14825 => x"20",
         14826 => x"70",
         14827 => x"62",
         14828 => x"66",
         14829 => x"73",
         14830 => x"65",
         14831 => x"6f",
         14832 => x"20",
         14833 => x"64",
         14834 => x"2e",
         14835 => x"73",
         14836 => x"6f",
         14837 => x"6e",
         14838 => x"65",
         14839 => x"00",
         14840 => x"69",
         14841 => x"6e",
         14842 => x"65",
         14843 => x"73",
         14844 => x"76",
         14845 => x"64",
         14846 => x"00",
         14847 => x"20",
         14848 => x"77",
         14849 => x"65",
         14850 => x"6f",
         14851 => x"74",
         14852 => x"00",
         14853 => x"6c",
         14854 => x"61",
         14855 => x"65",
         14856 => x"76",
         14857 => x"64",
         14858 => x"00",
         14859 => x"6c",
         14860 => x"6c",
         14861 => x"64",
         14862 => x"78",
         14863 => x"73",
         14864 => x"00",
         14865 => x"63",
         14866 => x"20",
         14867 => x"69",
         14868 => x"00",
         14869 => x"76",
         14870 => x"64",
         14871 => x"6c",
         14872 => x"6d",
         14873 => x"00",
         14874 => x"20",
         14875 => x"68",
         14876 => x"75",
         14877 => x"00",
         14878 => x"20",
         14879 => x"65",
         14880 => x"75",
         14881 => x"00",
         14882 => x"73",
         14883 => x"6f",
         14884 => x"65",
         14885 => x"2e",
         14886 => x"74",
         14887 => x"61",
         14888 => x"72",
         14889 => x"2e",
         14890 => x"73",
         14891 => x"72",
         14892 => x"00",
         14893 => x"63",
         14894 => x"73",
         14895 => x"00",
         14896 => x"6c",
         14897 => x"79",
         14898 => x"20",
         14899 => x"61",
         14900 => x"6c",
         14901 => x"79",
         14902 => x"2f",
         14903 => x"2e",
         14904 => x"00",
         14905 => x"61",
         14906 => x"00",
         14907 => x"38",
         14908 => x"00",
         14909 => x"20",
         14910 => x"32",
         14911 => x"00",
         14912 => x"00",
         14913 => x"00",
         14914 => x"00",
         14915 => x"34",
         14916 => x"00",
         14917 => x"20",
         14918 => x"20",
         14919 => x"00",
         14920 => x"53",
         14921 => x"20",
         14922 => x"28",
         14923 => x"2f",
         14924 => x"32",
         14925 => x"00",
         14926 => x"2e",
         14927 => x"00",
         14928 => x"50",
         14929 => x"72",
         14930 => x"25",
         14931 => x"29",
         14932 => x"20",
         14933 => x"2a",
         14934 => x"00",
         14935 => x"55",
         14936 => x"74",
         14937 => x"75",
         14938 => x"48",
         14939 => x"6c",
         14940 => x"00",
         14941 => x"52",
         14942 => x"54",
         14943 => x"6e",
         14944 => x"72",
         14945 => x"00",
         14946 => x"52",
         14947 => x"52",
         14948 => x"6e",
         14949 => x"72",
         14950 => x"00",
         14951 => x"52",
         14952 => x"54",
         14953 => x"6e",
         14954 => x"72",
         14955 => x"00",
         14956 => x"52",
         14957 => x"52",
         14958 => x"6e",
         14959 => x"72",
         14960 => x"00",
         14961 => x"43",
         14962 => x"57",
         14963 => x"6e",
         14964 => x"72",
         14965 => x"00",
         14966 => x"43",
         14967 => x"52",
         14968 => x"6e",
         14969 => x"72",
         14970 => x"00",
         14971 => x"32",
         14972 => x"74",
         14973 => x"75",
         14974 => x"00",
         14975 => x"6d",
         14976 => x"69",
         14977 => x"72",
         14978 => x"74",
         14979 => x"74",
         14980 => x"67",
         14981 => x"20",
         14982 => x"65",
         14983 => x"2e",
         14984 => x"61",
         14985 => x"6e",
         14986 => x"69",
         14987 => x"2e",
         14988 => x"00",
         14989 => x"74",
         14990 => x"65",
         14991 => x"61",
         14992 => x"00",
         14993 => x"53",
         14994 => x"75",
         14995 => x"74",
         14996 => x"69",
         14997 => x"20",
         14998 => x"69",
         14999 => x"69",
         15000 => x"73",
         15001 => x"64",
         15002 => x"72",
         15003 => x"2c",
         15004 => x"65",
         15005 => x"20",
         15006 => x"74",
         15007 => x"6e",
         15008 => x"6c",
         15009 => x"00",
         15010 => x"00",
         15011 => x"3a",
         15012 => x"00",
         15013 => x"00",
         15014 => x"64",
         15015 => x"6d",
         15016 => x"64",
         15017 => x"00",
         15018 => x"55",
         15019 => x"6e",
         15020 => x"3a",
         15021 => x"5c",
         15022 => x"25",
         15023 => x"00",
         15024 => x"6c",
         15025 => x"65",
         15026 => x"74",
         15027 => x"2e",
         15028 => x"00",
         15029 => x"73",
         15030 => x"74",
         15031 => x"20",
         15032 => x"6c",
         15033 => x"74",
         15034 => x"2e",
         15035 => x"00",
         15036 => x"6c",
         15037 => x"67",
         15038 => x"64",
         15039 => x"20",
         15040 => x"6c",
         15041 => x"2e",
         15042 => x"00",
         15043 => x"6c",
         15044 => x"65",
         15045 => x"6e",
         15046 => x"63",
         15047 => x"20",
         15048 => x"29",
         15049 => x"00",
         15050 => x"65",
         15051 => x"69",
         15052 => x"63",
         15053 => x"20",
         15054 => x"30",
         15055 => x"20",
         15056 => x"0a",
         15057 => x"38",
         15058 => x"25",
         15059 => x"58",
         15060 => x"00",
         15061 => x"38",
         15062 => x"25",
         15063 => x"2d",
         15064 => x"6d",
         15065 => x"69",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"38",
         15069 => x"25",
         15070 => x"29",
         15071 => x"30",
         15072 => x"28",
         15073 => x"78",
         15074 => x"00",
         15075 => x"70",
         15076 => x"67",
         15077 => x"00",
         15078 => x"38",
         15079 => x"25",
         15080 => x"2d",
         15081 => x"65",
         15082 => x"6e",
         15083 => x"2e",
         15084 => x"00",
         15085 => x"6d",
         15086 => x"65",
         15087 => x"79",
         15088 => x"6f",
         15089 => x"65",
         15090 => x"00",
         15091 => x"3a",
         15092 => x"5c",
         15093 => x"00",
         15094 => x"6d",
         15095 => x"20",
         15096 => x"61",
         15097 => x"65",
         15098 => x"63",
         15099 => x"6f",
         15100 => x"72",
         15101 => x"73",
         15102 => x"6f",
         15103 => x"6e",
         15104 => x"00",
         15105 => x"3f",
         15106 => x"2f",
         15107 => x"25",
         15108 => x"64",
         15109 => x"3a",
         15110 => x"25",
         15111 => x"0a",
         15112 => x"43",
         15113 => x"6e",
         15114 => x"75",
         15115 => x"69",
         15116 => x"00",
         15117 => x"44",
         15118 => x"63",
         15119 => x"69",
         15120 => x"65",
         15121 => x"74",
         15122 => x"00",
         15123 => x"64",
         15124 => x"73",
         15125 => x"00",
         15126 => x"20",
         15127 => x"55",
         15128 => x"73",
         15129 => x"56",
         15130 => x"6f",
         15131 => x"64",
         15132 => x"73",
         15133 => x"20",
         15134 => x"58",
         15135 => x"00",
         15136 => x"20",
         15137 => x"55",
         15138 => x"6d",
         15139 => x"20",
         15140 => x"72",
         15141 => x"64",
         15142 => x"73",
         15143 => x"20",
         15144 => x"58",
         15145 => x"00",
         15146 => x"20",
         15147 => x"61",
         15148 => x"53",
         15149 => x"74",
         15150 => x"64",
         15151 => x"73",
         15152 => x"20",
         15153 => x"20",
         15154 => x"58",
         15155 => x"00",
         15156 => x"73",
         15157 => x"00",
         15158 => x"20",
         15159 => x"55",
         15160 => x"20",
         15161 => x"20",
         15162 => x"20",
         15163 => x"20",
         15164 => x"20",
         15165 => x"20",
         15166 => x"58",
         15167 => x"00",
         15168 => x"20",
         15169 => x"73",
         15170 => x"20",
         15171 => x"63",
         15172 => x"72",
         15173 => x"20",
         15174 => x"20",
         15175 => x"20",
         15176 => x"25",
         15177 => x"4d",
         15178 => x"00",
         15179 => x"20",
         15180 => x"73",
         15181 => x"6e",
         15182 => x"44",
         15183 => x"20",
         15184 => x"63",
         15185 => x"72",
         15186 => x"20",
         15187 => x"25",
         15188 => x"4d",
         15189 => x"00",
         15190 => x"20",
         15191 => x"52",
         15192 => x"43",
         15193 => x"6b",
         15194 => x"65",
         15195 => x"20",
         15196 => x"20",
         15197 => x"20",
         15198 => x"25",
         15199 => x"4d",
         15200 => x"00",
         15201 => x"20",
         15202 => x"49",
         15203 => x"20",
         15204 => x"32",
         15205 => x"20",
         15206 => x"43",
         15207 => x"00",
         15208 => x"20",
         15209 => x"20",
         15210 => x"00",
         15211 => x"20",
         15212 => x"53",
         15213 => x"4e",
         15214 => x"55",
         15215 => x"00",
         15216 => x"20",
         15217 => x"54",
         15218 => x"54",
         15219 => x"28",
         15220 => x"6e",
         15221 => x"73",
         15222 => x"32",
         15223 => x"0a",
         15224 => x"20",
         15225 => x"4d",
         15226 => x"20",
         15227 => x"28",
         15228 => x"65",
         15229 => x"20",
         15230 => x"32",
         15231 => x"0a",
         15232 => x"20",
         15233 => x"20",
         15234 => x"44",
         15235 => x"28",
         15236 => x"69",
         15237 => x"20",
         15238 => x"32",
         15239 => x"0a",
         15240 => x"20",
         15241 => x"4d",
         15242 => x"20",
         15243 => x"28",
         15244 => x"58",
         15245 => x"38",
         15246 => x"0a",
         15247 => x"20",
         15248 => x"41",
         15249 => x"20",
         15250 => x"28",
         15251 => x"58",
         15252 => x"38",
         15253 => x"0a",
         15254 => x"20",
         15255 => x"53",
         15256 => x"52",
         15257 => x"28",
         15258 => x"58",
         15259 => x"38",
         15260 => x"0a",
         15261 => x"20",
         15262 => x"52",
         15263 => x"20",
         15264 => x"28",
         15265 => x"58",
         15266 => x"38",
         15267 => x"0a",
         15268 => x"20",
         15269 => x"20",
         15270 => x"41",
         15271 => x"28",
         15272 => x"58",
         15273 => x"38",
         15274 => x"0a",
         15275 => x"66",
         15276 => x"20",
         15277 => x"20",
         15278 => x"66",
         15279 => x"00",
         15280 => x"6b",
         15281 => x"6e",
         15282 => x"4f",
         15283 => x"00",
         15284 => x"61",
         15285 => x"00",
         15286 => x"64",
         15287 => x"00",
         15288 => x"65",
         15289 => x"00",
         15290 => x"4f",
         15291 => x"f0",
         15292 => x"00",
         15293 => x"00",
         15294 => x"f0",
         15295 => x"00",
         15296 => x"00",
         15297 => x"f0",
         15298 => x"00",
         15299 => x"00",
         15300 => x"f0",
         15301 => x"00",
         15302 => x"00",
         15303 => x"f0",
         15304 => x"00",
         15305 => x"00",
         15306 => x"f0",
         15307 => x"00",
         15308 => x"00",
         15309 => x"f0",
         15310 => x"00",
         15311 => x"00",
         15312 => x"f0",
         15313 => x"00",
         15314 => x"00",
         15315 => x"f0",
         15316 => x"00",
         15317 => x"00",
         15318 => x"f0",
         15319 => x"00",
         15320 => x"00",
         15321 => x"f0",
         15322 => x"00",
         15323 => x"00",
         15324 => x"f0",
         15325 => x"00",
         15326 => x"00",
         15327 => x"f0",
         15328 => x"00",
         15329 => x"00",
         15330 => x"f0",
         15331 => x"00",
         15332 => x"00",
         15333 => x"f0",
         15334 => x"00",
         15335 => x"00",
         15336 => x"f0",
         15337 => x"00",
         15338 => x"00",
         15339 => x"f0",
         15340 => x"00",
         15341 => x"00",
         15342 => x"f0",
         15343 => x"00",
         15344 => x"00",
         15345 => x"f0",
         15346 => x"00",
         15347 => x"00",
         15348 => x"ef",
         15349 => x"00",
         15350 => x"00",
         15351 => x"ef",
         15352 => x"00",
         15353 => x"00",
         15354 => x"ef",
         15355 => x"00",
         15356 => x"00",
         15357 => x"44",
         15358 => x"43",
         15359 => x"42",
         15360 => x"41",
         15361 => x"36",
         15362 => x"35",
         15363 => x"34",
         15364 => x"46",
         15365 => x"33",
         15366 => x"32",
         15367 => x"31",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"6e",
         15380 => x"20",
         15381 => x"6e",
         15382 => x"65",
         15383 => x"20",
         15384 => x"74",
         15385 => x"20",
         15386 => x"65",
         15387 => x"69",
         15388 => x"6c",
         15389 => x"2e",
         15390 => x"73",
         15391 => x"79",
         15392 => x"73",
         15393 => x"00",
         15394 => x"00",
         15395 => x"36",
         15396 => x"20",
         15397 => x"00",
         15398 => x"69",
         15399 => x"20",
         15400 => x"72",
         15401 => x"74",
         15402 => x"65",
         15403 => x"73",
         15404 => x"79",
         15405 => x"6c",
         15406 => x"6f",
         15407 => x"46",
         15408 => x"00",
         15409 => x"73",
         15410 => x"00",
         15411 => x"31",
         15412 => x"00",
         15413 => x"41",
         15414 => x"42",
         15415 => x"43",
         15416 => x"44",
         15417 => x"31",
         15418 => x"00",
         15419 => x"31",
         15420 => x"00",
         15421 => x"31",
         15422 => x"00",
         15423 => x"31",
         15424 => x"00",
         15425 => x"31",
         15426 => x"00",
         15427 => x"31",
         15428 => x"00",
         15429 => x"31",
         15430 => x"00",
         15431 => x"31",
         15432 => x"00",
         15433 => x"31",
         15434 => x"00",
         15435 => x"32",
         15436 => x"00",
         15437 => x"32",
         15438 => x"00",
         15439 => x"33",
         15440 => x"00",
         15441 => x"46",
         15442 => x"35",
         15443 => x"00",
         15444 => x"36",
         15445 => x"00",
         15446 => x"25",
         15447 => x"64",
         15448 => x"2c",
         15449 => x"25",
         15450 => x"64",
         15451 => x"32",
         15452 => x"00",
         15453 => x"25",
         15454 => x"64",
         15455 => x"3a",
         15456 => x"25",
         15457 => x"64",
         15458 => x"3a",
         15459 => x"2c",
         15460 => x"25",
         15461 => x"00",
         15462 => x"32",
         15463 => x"00",
         15464 => x"5b",
         15465 => x"25",
         15466 => x"00",
         15467 => x"70",
         15468 => x"20",
         15469 => x"73",
         15470 => x"00",
         15471 => x"3a",
         15472 => x"78",
         15473 => x"32",
         15474 => x"00",
         15475 => x"3a",
         15476 => x"78",
         15477 => x"32",
         15478 => x"00",
         15479 => x"3a",
         15480 => x"78",
         15481 => x"00",
         15482 => x"20",
         15483 => x"74",
         15484 => x"66",
         15485 => x"64",
         15486 => x"00",
         15487 => x"00",
         15488 => x"3a",
         15489 => x"7c",
         15490 => x"00",
         15491 => x"3b",
         15492 => x"00",
         15493 => x"54",
         15494 => x"54",
         15495 => x"00",
         15496 => x"90",
         15497 => x"4f",
         15498 => x"30",
         15499 => x"20",
         15500 => x"45",
         15501 => x"20",
         15502 => x"20",
         15503 => x"20",
         15504 => x"20",
         15505 => x"45",
         15506 => x"20",
         15507 => x"33",
         15508 => x"20",
         15509 => x"f1",
         15510 => x"00",
         15511 => x"00",
         15512 => x"00",
         15513 => x"05",
         15514 => x"10",
         15515 => x"18",
         15516 => x"00",
         15517 => x"45",
         15518 => x"8f",
         15519 => x"45",
         15520 => x"8e",
         15521 => x"92",
         15522 => x"55",
         15523 => x"9a",
         15524 => x"9e",
         15525 => x"4f",
         15526 => x"a6",
         15527 => x"aa",
         15528 => x"ae",
         15529 => x"b2",
         15530 => x"b6",
         15531 => x"ba",
         15532 => x"be",
         15533 => x"c2",
         15534 => x"c6",
         15535 => x"ca",
         15536 => x"ce",
         15537 => x"d2",
         15538 => x"d6",
         15539 => x"da",
         15540 => x"de",
         15541 => x"e2",
         15542 => x"e6",
         15543 => x"ea",
         15544 => x"ee",
         15545 => x"f2",
         15546 => x"f6",
         15547 => x"fa",
         15548 => x"fe",
         15549 => x"2c",
         15550 => x"5d",
         15551 => x"2a",
         15552 => x"3f",
         15553 => x"00",
         15554 => x"00",
         15555 => x"00",
         15556 => x"02",
         15557 => x"00",
         15558 => x"00",
         15559 => x"00",
         15560 => x"00",
         15561 => x"00",
         15562 => x"00",
         15563 => x"00",
         15564 => x"00",
         15565 => x"00",
         15566 => x"00",
         15567 => x"00",
         15568 => x"00",
         15569 => x"00",
         15570 => x"00",
         15571 => x"00",
         15572 => x"00",
         15573 => x"00",
         15574 => x"00",
         15575 => x"00",
         15576 => x"00",
         15577 => x"01",
         15578 => x"00",
         15579 => x"00",
         15580 => x"00",
         15581 => x"00",
         15582 => x"23",
         15583 => x"00",
         15584 => x"00",
         15585 => x"00",
         15586 => x"25",
         15587 => x"25",
         15588 => x"25",
         15589 => x"25",
         15590 => x"25",
         15591 => x"25",
         15592 => x"25",
         15593 => x"25",
         15594 => x"25",
         15595 => x"25",
         15596 => x"25",
         15597 => x"25",
         15598 => x"25",
         15599 => x"25",
         15600 => x"25",
         15601 => x"25",
         15602 => x"25",
         15603 => x"25",
         15604 => x"25",
         15605 => x"25",
         15606 => x"25",
         15607 => x"25",
         15608 => x"25",
         15609 => x"25",
         15610 => x"00",
         15611 => x"03",
         15612 => x"03",
         15613 => x"03",
         15614 => x"03",
         15615 => x"03",
         15616 => x"03",
         15617 => x"22",
         15618 => x"00",
         15619 => x"22",
         15620 => x"23",
         15621 => x"22",
         15622 => x"22",
         15623 => x"22",
         15624 => x"00",
         15625 => x"00",
         15626 => x"03",
         15627 => x"03",
         15628 => x"03",
         15629 => x"00",
         15630 => x"01",
         15631 => x"01",
         15632 => x"01",
         15633 => x"01",
         15634 => x"01",
         15635 => x"01",
         15636 => x"02",
         15637 => x"01",
         15638 => x"01",
         15639 => x"01",
         15640 => x"01",
         15641 => x"01",
         15642 => x"01",
         15643 => x"01",
         15644 => x"01",
         15645 => x"01",
         15646 => x"01",
         15647 => x"01",
         15648 => x"01",
         15649 => x"02",
         15650 => x"01",
         15651 => x"02",
         15652 => x"01",
         15653 => x"01",
         15654 => x"01",
         15655 => x"01",
         15656 => x"01",
         15657 => x"01",
         15658 => x"01",
         15659 => x"01",
         15660 => x"01",
         15661 => x"01",
         15662 => x"01",
         15663 => x"01",
         15664 => x"01",
         15665 => x"01",
         15666 => x"01",
         15667 => x"01",
         15668 => x"01",
         15669 => x"01",
         15670 => x"01",
         15671 => x"01",
         15672 => x"01",
         15673 => x"01",
         15674 => x"01",
         15675 => x"01",
         15676 => x"00",
         15677 => x"01",
         15678 => x"01",
         15679 => x"01",
         15680 => x"01",
         15681 => x"01",
         15682 => x"01",
         15683 => x"00",
         15684 => x"02",
         15685 => x"02",
         15686 => x"02",
         15687 => x"02",
         15688 => x"02",
         15689 => x"02",
         15690 => x"01",
         15691 => x"02",
         15692 => x"01",
         15693 => x"01",
         15694 => x"01",
         15695 => x"02",
         15696 => x"02",
         15697 => x"02",
         15698 => x"01",
         15699 => x"02",
         15700 => x"02",
         15701 => x"01",
         15702 => x"2c",
         15703 => x"02",
         15704 => x"01",
         15705 => x"02",
         15706 => x"02",
         15707 => x"01",
         15708 => x"02",
         15709 => x"02",
         15710 => x"02",
         15711 => x"2c",
         15712 => x"02",
         15713 => x"02",
         15714 => x"01",
         15715 => x"02",
         15716 => x"02",
         15717 => x"02",
         15718 => x"01",
         15719 => x"02",
         15720 => x"02",
         15721 => x"02",
         15722 => x"03",
         15723 => x"03",
         15724 => x"03",
         15725 => x"00",
         15726 => x"03",
         15727 => x"03",
         15728 => x"03",
         15729 => x"00",
         15730 => x"03",
         15731 => x"03",
         15732 => x"00",
         15733 => x"03",
         15734 => x"03",
         15735 => x"03",
         15736 => x"03",
         15737 => x"03",
         15738 => x"03",
         15739 => x"03",
         15740 => x"03",
         15741 => x"04",
         15742 => x"04",
         15743 => x"04",
         15744 => x"04",
         15745 => x"04",
         15746 => x"04",
         15747 => x"04",
         15748 => x"01",
         15749 => x"04",
         15750 => x"00",
         15751 => x"00",
         15752 => x"1e",
         15753 => x"1e",
         15754 => x"1f",
         15755 => x"1f",
         15756 => x"1f",
         15757 => x"1f",
         15758 => x"1f",
         15759 => x"1f",
         15760 => x"1f",
         15761 => x"1f",
         15762 => x"1f",
         15763 => x"1f",
         15764 => x"06",
         15765 => x"00",
         15766 => x"1f",
         15767 => x"1f",
         15768 => x"1f",
         15769 => x"1f",
         15770 => x"1f",
         15771 => x"1f",
         15772 => x"1f",
         15773 => x"06",
         15774 => x"06",
         15775 => x"06",
         15776 => x"00",
         15777 => x"1f",
         15778 => x"1f",
         15779 => x"00",
         15780 => x"1f",
         15781 => x"1f",
         15782 => x"1f",
         15783 => x"1f",
         15784 => x"00",
         15785 => x"21",
         15786 => x"21",
         15787 => x"02",
         15788 => x"00",
         15789 => x"24",
         15790 => x"2c",
         15791 => x"2c",
         15792 => x"2c",
         15793 => x"2c",
         15794 => x"2c",
         15795 => x"2d",
         15796 => x"ff",
         15797 => x"00",
         15798 => x"00",
         15799 => x"e6",
         15800 => x"01",
         15801 => x"00",
         15802 => x"00",
         15803 => x"e6",
         15804 => x"01",
         15805 => x"00",
         15806 => x"00",
         15807 => x"e6",
         15808 => x"03",
         15809 => x"00",
         15810 => x"00",
         15811 => x"e6",
         15812 => x"03",
         15813 => x"00",
         15814 => x"00",
         15815 => x"e6",
         15816 => x"03",
         15817 => x"00",
         15818 => x"00",
         15819 => x"e6",
         15820 => x"04",
         15821 => x"00",
         15822 => x"00",
         15823 => x"e6",
         15824 => x"04",
         15825 => x"00",
         15826 => x"00",
         15827 => x"e6",
         15828 => x"04",
         15829 => x"00",
         15830 => x"00",
         15831 => x"e6",
         15832 => x"04",
         15833 => x"00",
         15834 => x"00",
         15835 => x"e6",
         15836 => x"04",
         15837 => x"00",
         15838 => x"00",
         15839 => x"e6",
         15840 => x"04",
         15841 => x"00",
         15842 => x"00",
         15843 => x"e6",
         15844 => x"04",
         15845 => x"00",
         15846 => x"00",
         15847 => x"e6",
         15848 => x"05",
         15849 => x"00",
         15850 => x"00",
         15851 => x"e6",
         15852 => x"05",
         15853 => x"00",
         15854 => x"00",
         15855 => x"e6",
         15856 => x"05",
         15857 => x"00",
         15858 => x"00",
         15859 => x"e6",
         15860 => x"05",
         15861 => x"00",
         15862 => x"00",
         15863 => x"e6",
         15864 => x"07",
         15865 => x"00",
         15866 => x"00",
         15867 => x"e6",
         15868 => x"07",
         15869 => x"00",
         15870 => x"00",
         15871 => x"e6",
         15872 => x"08",
         15873 => x"00",
         15874 => x"00",
         15875 => x"e6",
         15876 => x"08",
         15877 => x"00",
         15878 => x"00",
         15879 => x"e6",
         15880 => x"08",
         15881 => x"00",
         15882 => x"00",
         15883 => x"e6",
         15884 => x"08",
         15885 => x"00",
         15886 => x"00",
         15887 => x"e6",
         15888 => x"08",
         15889 => x"00",
         15890 => x"00",
         15891 => x"e6",
         15892 => x"08",
         15893 => x"00",
         15894 => x"00",
         15895 => x"e6",
         15896 => x"09",
         15897 => x"00",
         15898 => x"00",
         15899 => x"e6",
         15900 => x"09",
         15901 => x"00",
         15902 => x"00",
         15903 => x"e7",
         15904 => x"09",
         15905 => x"00",
         15906 => x"00",
         15907 => x"e7",
         15908 => x"09",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"7f",
         15914 => x"00",
         15915 => x"7f",
         15916 => x"00",
         15917 => x"7f",
         15918 => x"00",
         15919 => x"00",
         15920 => x"00",
         15921 => x"ff",
         15922 => x"00",
         15923 => x"00",
         15924 => x"78",
         15925 => x"00",
         15926 => x"e1",
         15927 => x"e1",
         15928 => x"e1",
         15929 => x"00",
         15930 => x"01",
         15931 => x"01",
         15932 => x"10",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"f0",
         15959 => x"00",
         15960 => x"f0",
         15961 => x"00",
         15962 => x"f0",
         15963 => x"00",
         15964 => x"fd",
         15965 => x"5f",
         15966 => x"3a",
         15967 => x"40",
         15968 => x"f0",
         15969 => x"73",
         15970 => x"77",
         15971 => x"6b",
         15972 => x"6f",
         15973 => x"63",
         15974 => x"67",
         15975 => x"33",
         15976 => x"37",
         15977 => x"2d",
         15978 => x"2c",
         15979 => x"f3",
         15980 => x"3f",
         15981 => x"f0",
         15982 => x"f0",
         15983 => x"82",
         15984 => x"f0",
         15985 => x"58",
         15986 => x"3b",
         15987 => x"40",
         15988 => x"f0",
         15989 => x"53",
         15990 => x"57",
         15991 => x"4b",
         15992 => x"4f",
         15993 => x"43",
         15994 => x"47",
         15995 => x"33",
         15996 => x"37",
         15997 => x"2d",
         15998 => x"2c",
         15999 => x"f3",
         16000 => x"3f",
         16001 => x"f0",
         16002 => x"f0",
         16003 => x"82",
         16004 => x"f0",
         16005 => x"58",
         16006 => x"2a",
         16007 => x"60",
         16008 => x"f0",
         16009 => x"53",
         16010 => x"57",
         16011 => x"4b",
         16012 => x"4f",
         16013 => x"43",
         16014 => x"47",
         16015 => x"23",
         16016 => x"27",
         16017 => x"3d",
         16018 => x"3c",
         16019 => x"e0",
         16020 => x"3f",
         16021 => x"f0",
         16022 => x"f0",
         16023 => x"87",
         16024 => x"f0",
         16025 => x"1e",
         16026 => x"f0",
         16027 => x"00",
         16028 => x"f0",
         16029 => x"13",
         16030 => x"17",
         16031 => x"0b",
         16032 => x"0f",
         16033 => x"03",
         16034 => x"07",
         16035 => x"f0",
         16036 => x"f0",
         16037 => x"f0",
         16038 => x"f0",
         16039 => x"f0",
         16040 => x"f0",
         16041 => x"f0",
         16042 => x"f0",
         16043 => x"82",
         16044 => x"f0",
         16045 => x"cf",
         16046 => x"4d",
         16047 => x"d7",
         16048 => x"f0",
         16049 => x"41",
         16050 => x"78",
         16051 => x"6c",
         16052 => x"d5",
         16053 => x"d9",
         16054 => x"4c",
         16055 => x"7e",
         16056 => x"5f",
         16057 => x"d1",
         16058 => x"d0",
         16059 => x"c2",
         16060 => x"bb",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"82",
         16064 => x"f0",
         16065 => x"00",
         16066 => x"00",
         16067 => x"00",
         16068 => x"00",
         16069 => x"00",
         16070 => x"00",
         16071 => x"00",
         16072 => x"00",
         16073 => x"00",
         16074 => x"00",
         16075 => x"00",
         16076 => x"00",
         16077 => x"00",
         16078 => x"00",
         16079 => x"00",
         16080 => x"00",
         16081 => x"00",
         16082 => x"00",
         16083 => x"00",
         16084 => x"00",
         16085 => x"00",
         16086 => x"00",
         16087 => x"00",
         16088 => x"00",
         16089 => x"00",
         16090 => x"00",
         16091 => x"00",
         16092 => x"00",
         16093 => x"f0",
         16094 => x"00",
         16095 => x"f0",
         16096 => x"00",
         16097 => x"f0",
         16098 => x"00",
         16099 => x"f0",
         16100 => x"00",
         16101 => x"f0",
         16102 => x"00",
         16103 => x"f0",
         16104 => x"00",
         16105 => x"f0",
         16106 => x"00",
         16107 => x"f0",
         16108 => x"00",
         16109 => x"f0",
         16110 => x"00",
         16111 => x"f1",
         16112 => x"00",
         16113 => x"f1",
         16114 => x"00",
         16115 => x"f1",
         16116 => x"00",
         16117 => x"f1",
         16118 => x"00",
         16119 => x"f1",
         16120 => x"00",
         16121 => x"f1",
         16122 => x"00",
         16123 => x"f1",
         16124 => x"00",
         16125 => x"f1",
         16126 => x"00",
         16127 => x"f1",
         16128 => x"00",
         16129 => x"f1",
         16130 => x"00",
         16131 => x"f1",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"32",
         18134 => x"01",
         18135 => x"00",
         18136 => x"f2",
         18137 => x"f6",
         18138 => x"fa",
         18139 => x"fe",
         18140 => x"c2",
         18141 => x"c6",
         18142 => x"e5",
         18143 => x"ef",
         18144 => x"62",
         18145 => x"66",
         18146 => x"6b",
         18147 => x"2e",
         18148 => x"22",
         18149 => x"26",
         18150 => x"4f",
         18151 => x"57",
         18152 => x"02",
         18153 => x"06",
         18154 => x"0a",
         18155 => x"0e",
         18156 => x"12",
         18157 => x"16",
         18158 => x"1a",
         18159 => x"be",
         18160 => x"82",
         18161 => x"86",
         18162 => x"8a",
         18163 => x"8e",
         18164 => x"92",
         18165 => x"96",
         18166 => x"9a",
         18167 => x"a5",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"01",
         18200 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"b5",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"91",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"92",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"84",
           386 => x"80",
           387 => x"84",
           388 => x"80",
           389 => x"04",
           390 => x"0c",
           391 => x"84",
           392 => x"80",
           393 => x"04",
           394 => x"0c",
           395 => x"84",
           396 => x"80",
           397 => x"04",
           398 => x"0c",
           399 => x"84",
           400 => x"80",
           401 => x"04",
           402 => x"0c",
           403 => x"84",
           404 => x"80",
           405 => x"04",
           406 => x"0c",
           407 => x"84",
           408 => x"80",
           409 => x"04",
           410 => x"0c",
           411 => x"84",
           412 => x"80",
           413 => x"04",
           414 => x"0c",
           415 => x"84",
           416 => x"80",
           417 => x"04",
           418 => x"0c",
           419 => x"84",
           420 => x"80",
           421 => x"04",
           422 => x"0c",
           423 => x"84",
           424 => x"80",
           425 => x"04",
           426 => x"0c",
           427 => x"84",
           428 => x"80",
           429 => x"04",
           430 => x"0c",
           431 => x"84",
           432 => x"80",
           433 => x"04",
           434 => x"0c",
           435 => x"2d",
           436 => x"08",
           437 => x"90",
           438 => x"f0",
           439 => x"b6",
           440 => x"f0",
           441 => x"80",
           442 => x"b8",
           443 => x"d2",
           444 => x"b8",
           445 => x"c0",
           446 => x"84",
           447 => x"80",
           448 => x"84",
           449 => x"80",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"90",
           455 => x"f0",
           456 => x"ef",
           457 => x"f0",
           458 => x"80",
           459 => x"b8",
           460 => x"d2",
           461 => x"b8",
           462 => x"c0",
           463 => x"84",
           464 => x"82",
           465 => x"84",
           466 => x"80",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"90",
           472 => x"f0",
           473 => x"94",
           474 => x"f0",
           475 => x"80",
           476 => x"b8",
           477 => x"de",
           478 => x"b8",
           479 => x"c0",
           480 => x"84",
           481 => x"82",
           482 => x"84",
           483 => x"80",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"90",
           489 => x"f0",
           490 => x"cf",
           491 => x"f0",
           492 => x"80",
           493 => x"b8",
           494 => x"84",
           495 => x"b8",
           496 => x"c0",
           497 => x"84",
           498 => x"82",
           499 => x"84",
           500 => x"80",
           501 => x"04",
           502 => x"0c",
           503 => x"2d",
           504 => x"08",
           505 => x"90",
           506 => x"f0",
           507 => x"ac",
           508 => x"f0",
           509 => x"80",
           510 => x"b8",
           511 => x"93",
           512 => x"b8",
           513 => x"c0",
           514 => x"84",
           515 => x"83",
           516 => x"84",
           517 => x"80",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"90",
           523 => x"f0",
           524 => x"d6",
           525 => x"f0",
           526 => x"80",
           527 => x"b8",
           528 => x"e6",
           529 => x"b8",
           530 => x"c0",
           531 => x"84",
           532 => x"82",
           533 => x"84",
           534 => x"80",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"90",
           540 => x"f0",
           541 => x"e6",
           542 => x"f0",
           543 => x"80",
           544 => x"b8",
           545 => x"a0",
           546 => x"b8",
           547 => x"c0",
           548 => x"84",
           549 => x"82",
           550 => x"84",
           551 => x"80",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"90",
           557 => x"f0",
           558 => x"82",
           559 => x"f0",
           560 => x"80",
           561 => x"b8",
           562 => x"b7",
           563 => x"b8",
           564 => x"c0",
           565 => x"84",
           566 => x"81",
           567 => x"84",
           568 => x"80",
           569 => x"04",
           570 => x"0c",
           571 => x"2d",
           572 => x"08",
           573 => x"90",
           574 => x"f0",
           575 => x"d0",
           576 => x"f0",
           577 => x"80",
           578 => x"b8",
           579 => x"d0",
           580 => x"b8",
           581 => x"c0",
           582 => x"84",
           583 => x"80",
           584 => x"84",
           585 => x"80",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"90",
           591 => x"f0",
           592 => x"2d",
           593 => x"08",
           594 => x"90",
           595 => x"f0",
           596 => x"f0",
           597 => x"f0",
           598 => x"80",
           599 => x"b8",
           600 => x"dc",
           601 => x"b8",
           602 => x"c0",
           603 => x"84",
           604 => x"81",
           605 => x"84",
           606 => x"80",
           607 => x"04",
           608 => x"0c",
           609 => x"2d",
           610 => x"08",
           611 => x"90",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"51",
           621 => x"73",
           622 => x"73",
           623 => x"81",
           624 => x"10",
           625 => x"07",
           626 => x"0c",
           627 => x"72",
           628 => x"81",
           629 => x"09",
           630 => x"71",
           631 => x"0a",
           632 => x"72",
           633 => x"51",
           634 => x"84",
           635 => x"84",
           636 => x"8e",
           637 => x"70",
           638 => x"0c",
           639 => x"93",
           640 => x"81",
           641 => x"ba",
           642 => x"3d",
           643 => x"70",
           644 => x"52",
           645 => x"74",
           646 => x"c8",
           647 => x"c5",
           648 => x"0d",
           649 => x"0d",
           650 => x"85",
           651 => x"32",
           652 => x"73",
           653 => x"58",
           654 => x"52",
           655 => x"09",
           656 => x"d3",
           657 => x"77",
           658 => x"70",
           659 => x"07",
           660 => x"55",
           661 => x"80",
           662 => x"38",
           663 => x"b2",
           664 => x"8e",
           665 => x"b8",
           666 => x"84",
           667 => x"ff",
           668 => x"84",
           669 => x"75",
           670 => x"57",
           671 => x"73",
           672 => x"30",
           673 => x"9f",
           674 => x"54",
           675 => x"24",
           676 => x"75",
           677 => x"71",
           678 => x"0c",
           679 => x"04",
           680 => x"b8",
           681 => x"3d",
           682 => x"3d",
           683 => x"86",
           684 => x"99",
           685 => x"56",
           686 => x"8e",
           687 => x"53",
           688 => x"3d",
           689 => x"9d",
           690 => x"54",
           691 => x"8d",
           692 => x"fd",
           693 => x"3d",
           694 => x"76",
           695 => x"85",
           696 => x"0d",
           697 => x"0d",
           698 => x"42",
           699 => x"70",
           700 => x"85",
           701 => x"81",
           702 => x"81",
           703 => x"5b",
           704 => x"7b",
           705 => x"06",
           706 => x"7b",
           707 => x"7b",
           708 => x"38",
           709 => x"81",
           710 => x"72",
           711 => x"81",
           712 => x"5f",
           713 => x"81",
           714 => x"b0",
           715 => x"70",
           716 => x"54",
           717 => x"38",
           718 => x"a9",
           719 => x"2a",
           720 => x"81",
           721 => x"7e",
           722 => x"38",
           723 => x"07",
           724 => x"57",
           725 => x"38",
           726 => x"54",
           727 => x"e4",
           728 => x"0d",
           729 => x"2a",
           730 => x"10",
           731 => x"05",
           732 => x"70",
           733 => x"70",
           734 => x"29",
           735 => x"70",
           736 => x"5a",
           737 => x"80",
           738 => x"86",
           739 => x"06",
           740 => x"bd",
           741 => x"33",
           742 => x"fe",
           743 => x"b8",
           744 => x"2e",
           745 => x"93",
           746 => x"74",
           747 => x"8a",
           748 => x"5a",
           749 => x"38",
           750 => x"7c",
           751 => x"8b",
           752 => x"33",
           753 => x"cc",
           754 => x"39",
           755 => x"70",
           756 => x"55",
           757 => x"81",
           758 => x"40",
           759 => x"38",
           760 => x"72",
           761 => x"97",
           762 => x"10",
           763 => x"05",
           764 => x"04",
           765 => x"54",
           766 => x"73",
           767 => x"7c",
           768 => x"8a",
           769 => x"7c",
           770 => x"76",
           771 => x"fe",
           772 => x"ff",
           773 => x"39",
           774 => x"60",
           775 => x"08",
           776 => x"cf",
           777 => x"41",
           778 => x"f4",
           779 => x"75",
           780 => x"3f",
           781 => x"08",
           782 => x"84",
           783 => x"18",
           784 => x"53",
           785 => x"88",
           786 => x"e4",
           787 => x"55",
           788 => x"81",
           789 => x"79",
           790 => x"90",
           791 => x"b8",
           792 => x"84",
           793 => x"c5",
           794 => x"b8",
           795 => x"2b",
           796 => x"40",
           797 => x"2e",
           798 => x"84",
           799 => x"fc",
           800 => x"70",
           801 => x"55",
           802 => x"70",
           803 => x"5f",
           804 => x"9e",
           805 => x"80",
           806 => x"80",
           807 => x"79",
           808 => x"38",
           809 => x"80",
           810 => x"80",
           811 => x"90",
           812 => x"83",
           813 => x"06",
           814 => x"80",
           815 => x"75",
           816 => x"81",
           817 => x"54",
           818 => x"86",
           819 => x"83",
           820 => x"70",
           821 => x"86",
           822 => x"5b",
           823 => x"54",
           824 => x"85",
           825 => x"79",
           826 => x"70",
           827 => x"83",
           828 => x"59",
           829 => x"2e",
           830 => x"7a",
           831 => x"06",
           832 => x"eb",
           833 => x"2a",
           834 => x"73",
           835 => x"7a",
           836 => x"06",
           837 => x"97",
           838 => x"06",
           839 => x"8f",
           840 => x"2a",
           841 => x"7e",
           842 => x"38",
           843 => x"80",
           844 => x"80",
           845 => x"90",
           846 => x"54",
           847 => x"9d",
           848 => x"b0",
           849 => x"3f",
           850 => x"80",
           851 => x"80",
           852 => x"90",
           853 => x"54",
           854 => x"e5",
           855 => x"06",
           856 => x"2e",
           857 => x"79",
           858 => x"29",
           859 => x"05",
           860 => x"5b",
           861 => x"75",
           862 => x"7c",
           863 => x"87",
           864 => x"79",
           865 => x"29",
           866 => x"05",
           867 => x"5b",
           868 => x"80",
           869 => x"7a",
           870 => x"81",
           871 => x"7a",
           872 => x"b9",
           873 => x"e3",
           874 => x"38",
           875 => x"2e",
           876 => x"76",
           877 => x"81",
           878 => x"84",
           879 => x"96",
           880 => x"ff",
           881 => x"52",
           882 => x"3f",
           883 => x"f4",
           884 => x"06",
           885 => x"81",
           886 => x"80",
           887 => x"38",
           888 => x"80",
           889 => x"80",
           890 => x"90",
           891 => x"55",
           892 => x"fc",
           893 => x"52",
           894 => x"f4",
           895 => x"7a",
           896 => x"7a",
           897 => x"33",
           898 => x"fa",
           899 => x"c8",
           900 => x"c0",
           901 => x"f8",
           902 => x"61",
           903 => x"08",
           904 => x"cf",
           905 => x"42",
           906 => x"fd",
           907 => x"84",
           908 => x"80",
           909 => x"13",
           910 => x"2b",
           911 => x"84",
           912 => x"fc",
           913 => x"70",
           914 => x"52",
           915 => x"41",
           916 => x"2a",
           917 => x"5c",
           918 => x"c9",
           919 => x"84",
           920 => x"fc",
           921 => x"70",
           922 => x"54",
           923 => x"25",
           924 => x"7c",
           925 => x"85",
           926 => x"39",
           927 => x"83",
           928 => x"5b",
           929 => x"ff",
           930 => x"ca",
           931 => x"75",
           932 => x"57",
           933 => x"d8",
           934 => x"ff",
           935 => x"ff",
           936 => x"54",
           937 => x"ff",
           938 => x"38",
           939 => x"70",
           940 => x"33",
           941 => x"3f",
           942 => x"fc",
           943 => x"fc",
           944 => x"84",
           945 => x"fc",
           946 => x"70",
           947 => x"58",
           948 => x"7b",
           949 => x"81",
           950 => x"57",
           951 => x"38",
           952 => x"7f",
           953 => x"71",
           954 => x"40",
           955 => x"7e",
           956 => x"38",
           957 => x"bf",
           958 => x"b8",
           959 => x"ad",
           960 => x"07",
           961 => x"5b",
           962 => x"38",
           963 => x"7a",
           964 => x"80",
           965 => x"59",
           966 => x"38",
           967 => x"7f",
           968 => x"71",
           969 => x"06",
           970 => x"5f",
           971 => x"38",
           972 => x"f6",
           973 => x"e4",
           974 => x"ff",
           975 => x"31",
           976 => x"5a",
           977 => x"58",
           978 => x"7a",
           979 => x"7c",
           980 => x"76",
           981 => x"f7",
           982 => x"60",
           983 => x"08",
           984 => x"5d",
           985 => x"79",
           986 => x"75",
           987 => x"3f",
           988 => x"08",
           989 => x"06",
           990 => x"90",
           991 => x"c4",
           992 => x"80",
           993 => x"58",
           994 => x"88",
           995 => x"39",
           996 => x"80",
           997 => x"80",
           998 => x"90",
           999 => x"54",
          1000 => x"fa",
          1001 => x"52",
          1002 => x"c4",
          1003 => x"7c",
          1004 => x"83",
          1005 => x"90",
          1006 => x"06",
          1007 => x"7c",
          1008 => x"83",
          1009 => x"88",
          1010 => x"5f",
          1011 => x"fb",
          1012 => x"d8",
          1013 => x"2c",
          1014 => x"90",
          1015 => x"2c",
          1016 => x"06",
          1017 => x"53",
          1018 => x"38",
          1019 => x"7c",
          1020 => x"82",
          1021 => x"81",
          1022 => x"80",
          1023 => x"38",
          1024 => x"7c",
          1025 => x"2a",
          1026 => x"3f",
          1027 => x"5b",
          1028 => x"f7",
          1029 => x"c8",
          1030 => x"31",
          1031 => x"98",
          1032 => x"f9",
          1033 => x"52",
          1034 => x"c4",
          1035 => x"7c",
          1036 => x"82",
          1037 => x"be",
          1038 => x"75",
          1039 => x"3f",
          1040 => x"08",
          1041 => x"06",
          1042 => x"90",
          1043 => x"fd",
          1044 => x"82",
          1045 => x"71",
          1046 => x"06",
          1047 => x"fd",
          1048 => x"3d",
          1049 => x"c4",
          1050 => x"52",
          1051 => x"b5",
          1052 => x"0d",
          1053 => x"0d",
          1054 => x"0b",
          1055 => x"08",
          1056 => x"70",
          1057 => x"32",
          1058 => x"51",
          1059 => x"57",
          1060 => x"77",
          1061 => x"06",
          1062 => x"74",
          1063 => x"56",
          1064 => x"77",
          1065 => x"84",
          1066 => x"52",
          1067 => x"14",
          1068 => x"2d",
          1069 => x"08",
          1070 => x"38",
          1071 => x"70",
          1072 => x"33",
          1073 => x"2e",
          1074 => x"d4",
          1075 => x"d7",
          1076 => x"c8",
          1077 => x"d4",
          1078 => x"8a",
          1079 => x"08",
          1080 => x"84",
          1081 => x"80",
          1082 => x"ff",
          1083 => x"75",
          1084 => x"0c",
          1085 => x"04",
          1086 => x"78",
          1087 => x"80",
          1088 => x"33",
          1089 => x"81",
          1090 => x"06",
          1091 => x"57",
          1092 => x"77",
          1093 => x"06",
          1094 => x"70",
          1095 => x"33",
          1096 => x"2e",
          1097 => x"98",
          1098 => x"75",
          1099 => x"0c",
          1100 => x"04",
          1101 => x"05",
          1102 => x"72",
          1103 => x"38",
          1104 => x"51",
          1105 => x"53",
          1106 => x"b8",
          1107 => x"2e",
          1108 => x"74",
          1109 => x"56",
          1110 => x"72",
          1111 => x"39",
          1112 => x"84",
          1113 => x"52",
          1114 => x"3f",
          1115 => x"04",
          1116 => x"78",
          1117 => x"33",
          1118 => x"81",
          1119 => x"56",
          1120 => x"ff",
          1121 => x"38",
          1122 => x"81",
          1123 => x"80",
          1124 => x"8c",
          1125 => x"72",
          1126 => x"25",
          1127 => x"08",
          1128 => x"34",
          1129 => x"05",
          1130 => x"15",
          1131 => x"13",
          1132 => x"76",
          1133 => x"b8",
          1134 => x"3d",
          1135 => x"52",
          1136 => x"06",
          1137 => x"08",
          1138 => x"ff",
          1139 => x"e4",
          1140 => x"8c",
          1141 => x"05",
          1142 => x"76",
          1143 => x"fb",
          1144 => x"85",
          1145 => x"81",
          1146 => x"81",
          1147 => x"55",
          1148 => x"ff",
          1149 => x"38",
          1150 => x"81",
          1151 => x"b3",
          1152 => x"2a",
          1153 => x"71",
          1154 => x"c3",
          1155 => x"70",
          1156 => x"71",
          1157 => x"f0",
          1158 => x"76",
          1159 => x"08",
          1160 => x"17",
          1161 => x"ff",
          1162 => x"84",
          1163 => x"87",
          1164 => x"74",
          1165 => x"53",
          1166 => x"34",
          1167 => x"81",
          1168 => x"0c",
          1169 => x"84",
          1170 => x"87",
          1171 => x"75",
          1172 => x"08",
          1173 => x"84",
          1174 => x"52",
          1175 => x"08",
          1176 => x"b9",
          1177 => x"33",
          1178 => x"54",
          1179 => x"e4",
          1180 => x"85",
          1181 => x"07",
          1182 => x"17",
          1183 => x"73",
          1184 => x"0c",
          1185 => x"04",
          1186 => x"53",
          1187 => x"34",
          1188 => x"39",
          1189 => x"75",
          1190 => x"54",
          1191 => x"81",
          1192 => x"51",
          1193 => x"ff",
          1194 => x"70",
          1195 => x"33",
          1196 => x"70",
          1197 => x"34",
          1198 => x"73",
          1199 => x"0c",
          1200 => x"04",
          1201 => x"76",
          1202 => x"55",
          1203 => x"70",
          1204 => x"38",
          1205 => x"a1",
          1206 => x"2e",
          1207 => x"70",
          1208 => x"33",
          1209 => x"05",
          1210 => x"11",
          1211 => x"38",
          1212 => x"e4",
          1213 => x"0d",
          1214 => x"55",
          1215 => x"d9",
          1216 => x"75",
          1217 => x"13",
          1218 => x"53",
          1219 => x"34",
          1220 => x"70",
          1221 => x"38",
          1222 => x"13",
          1223 => x"33",
          1224 => x"11",
          1225 => x"38",
          1226 => x"3d",
          1227 => x"53",
          1228 => x"81",
          1229 => x"51",
          1230 => x"ff",
          1231 => x"31",
          1232 => x"0c",
          1233 => x"0d",
          1234 => x"0d",
          1235 => x"54",
          1236 => x"70",
          1237 => x"33",
          1238 => x"70",
          1239 => x"34",
          1240 => x"73",
          1241 => x"0c",
          1242 => x"04",
          1243 => x"75",
          1244 => x"55",
          1245 => x"70",
          1246 => x"38",
          1247 => x"05",
          1248 => x"70",
          1249 => x"34",
          1250 => x"70",
          1251 => x"84",
          1252 => x"85",
          1253 => x"fc",
          1254 => x"78",
          1255 => x"54",
          1256 => x"a1",
          1257 => x"75",
          1258 => x"57",
          1259 => x"71",
          1260 => x"81",
          1261 => x"81",
          1262 => x"80",
          1263 => x"ff",
          1264 => x"e1",
          1265 => x"70",
          1266 => x"0c",
          1267 => x"04",
          1268 => x"f1",
          1269 => x"53",
          1270 => x"80",
          1271 => x"ff",
          1272 => x"81",
          1273 => x"2e",
          1274 => x"72",
          1275 => x"e4",
          1276 => x"0d",
          1277 => x"b8",
          1278 => x"3d",
          1279 => x"3d",
          1280 => x"53",
          1281 => x"80",
          1282 => x"b8",
          1283 => x"b8",
          1284 => x"05",
          1285 => x"b2",
          1286 => x"b8",
          1287 => x"84",
          1288 => x"80",
          1289 => x"84",
          1290 => x"15",
          1291 => x"34",
          1292 => x"52",
          1293 => x"08",
          1294 => x"3f",
          1295 => x"08",
          1296 => x"b8",
          1297 => x"3d",
          1298 => x"3d",
          1299 => x"71",
          1300 => x"53",
          1301 => x"2e",
          1302 => x"70",
          1303 => x"33",
          1304 => x"2e",
          1305 => x"12",
          1306 => x"2e",
          1307 => x"ea",
          1308 => x"70",
          1309 => x"52",
          1310 => x"e4",
          1311 => x"0d",
          1312 => x"0d",
          1313 => x"72",
          1314 => x"54",
          1315 => x"8e",
          1316 => x"70",
          1317 => x"34",
          1318 => x"70",
          1319 => x"84",
          1320 => x"85",
          1321 => x"fa",
          1322 => x"7a",
          1323 => x"52",
          1324 => x"8b",
          1325 => x"80",
          1326 => x"b8",
          1327 => x"e0",
          1328 => x"80",
          1329 => x"73",
          1330 => x"3f",
          1331 => x"e4",
          1332 => x"80",
          1333 => x"26",
          1334 => x"73",
          1335 => x"2e",
          1336 => x"81",
          1337 => x"2a",
          1338 => x"76",
          1339 => x"54",
          1340 => x"56",
          1341 => x"a8",
          1342 => x"74",
          1343 => x"74",
          1344 => x"78",
          1345 => x"11",
          1346 => x"81",
          1347 => x"06",
          1348 => x"ff",
          1349 => x"52",
          1350 => x"55",
          1351 => x"38",
          1352 => x"07",
          1353 => x"b8",
          1354 => x"3d",
          1355 => x"3d",
          1356 => x"fc",
          1357 => x"70",
          1358 => x"07",
          1359 => x"84",
          1360 => x"31",
          1361 => x"70",
          1362 => x"06",
          1363 => x"80",
          1364 => x"88",
          1365 => x"71",
          1366 => x"f0",
          1367 => x"70",
          1368 => x"2b",
          1369 => x"74",
          1370 => x"53",
          1371 => x"73",
          1372 => x"30",
          1373 => x"10",
          1374 => x"77",
          1375 => x"81",
          1376 => x"70",
          1377 => x"30",
          1378 => x"06",
          1379 => x"84",
          1380 => x"51",
          1381 => x"51",
          1382 => x"53",
          1383 => x"51",
          1384 => x"56",
          1385 => x"54",
          1386 => x"0d",
          1387 => x"0d",
          1388 => x"54",
          1389 => x"54",
          1390 => x"84",
          1391 => x"73",
          1392 => x"31",
          1393 => x"0c",
          1394 => x"0d",
          1395 => x"0d",
          1396 => x"54",
          1397 => x"80",
          1398 => x"76",
          1399 => x"3f",
          1400 => x"08",
          1401 => x"52",
          1402 => x"8d",
          1403 => x"fe",
          1404 => x"84",
          1405 => x"31",
          1406 => x"71",
          1407 => x"c5",
          1408 => x"71",
          1409 => x"38",
          1410 => x"71",
          1411 => x"31",
          1412 => x"57",
          1413 => x"80",
          1414 => x"2e",
          1415 => x"10",
          1416 => x"07",
          1417 => x"07",
          1418 => x"ff",
          1419 => x"70",
          1420 => x"72",
          1421 => x"31",
          1422 => x"56",
          1423 => x"58",
          1424 => x"da",
          1425 => x"b8",
          1426 => x"3d",
          1427 => x"3d",
          1428 => x"2c",
          1429 => x"7a",
          1430 => x"32",
          1431 => x"7d",
          1432 => x"32",
          1433 => x"57",
          1434 => x"56",
          1435 => x"55",
          1436 => x"3f",
          1437 => x"08",
          1438 => x"31",
          1439 => x"0c",
          1440 => x"04",
          1441 => x"7b",
          1442 => x"80",
          1443 => x"77",
          1444 => x"56",
          1445 => x"a0",
          1446 => x"06",
          1447 => x"15",
          1448 => x"70",
          1449 => x"73",
          1450 => x"38",
          1451 => x"80",
          1452 => x"b0",
          1453 => x"38",
          1454 => x"80",
          1455 => x"26",
          1456 => x"8a",
          1457 => x"a0",
          1458 => x"c4",
          1459 => x"74",
          1460 => x"e0",
          1461 => x"ff",
          1462 => x"d0",
          1463 => x"ff",
          1464 => x"90",
          1465 => x"38",
          1466 => x"81",
          1467 => x"54",
          1468 => x"81",
          1469 => x"78",
          1470 => x"38",
          1471 => x"13",
          1472 => x"79",
          1473 => x"56",
          1474 => x"a0",
          1475 => x"38",
          1476 => x"84",
          1477 => x"56",
          1478 => x"81",
          1479 => x"b8",
          1480 => x"3d",
          1481 => x"70",
          1482 => x"0c",
          1483 => x"56",
          1484 => x"2e",
          1485 => x"fe",
          1486 => x"15",
          1487 => x"70",
          1488 => x"73",
          1489 => x"a6",
          1490 => x"73",
          1491 => x"a0",
          1492 => x"a0",
          1493 => x"38",
          1494 => x"80",
          1495 => x"89",
          1496 => x"e1",
          1497 => x"b8",
          1498 => x"3d",
          1499 => x"58",
          1500 => x"78",
          1501 => x"55",
          1502 => x"fe",
          1503 => x"0b",
          1504 => x"0c",
          1505 => x"04",
          1506 => x"7b",
          1507 => x"80",
          1508 => x"77",
          1509 => x"56",
          1510 => x"a0",
          1511 => x"06",
          1512 => x"15",
          1513 => x"70",
          1514 => x"73",
          1515 => x"38",
          1516 => x"80",
          1517 => x"b0",
          1518 => x"38",
          1519 => x"80",
          1520 => x"26",
          1521 => x"8a",
          1522 => x"a0",
          1523 => x"c4",
          1524 => x"74",
          1525 => x"e0",
          1526 => x"ff",
          1527 => x"d0",
          1528 => x"ff",
          1529 => x"90",
          1530 => x"38",
          1531 => x"81",
          1532 => x"54",
          1533 => x"81",
          1534 => x"78",
          1535 => x"38",
          1536 => x"13",
          1537 => x"79",
          1538 => x"56",
          1539 => x"a0",
          1540 => x"38",
          1541 => x"84",
          1542 => x"56",
          1543 => x"81",
          1544 => x"b8",
          1545 => x"3d",
          1546 => x"70",
          1547 => x"0c",
          1548 => x"56",
          1549 => x"2e",
          1550 => x"fe",
          1551 => x"15",
          1552 => x"70",
          1553 => x"73",
          1554 => x"a6",
          1555 => x"73",
          1556 => x"a0",
          1557 => x"a0",
          1558 => x"38",
          1559 => x"80",
          1560 => x"89",
          1561 => x"e1",
          1562 => x"b8",
          1563 => x"3d",
          1564 => x"58",
          1565 => x"78",
          1566 => x"55",
          1567 => x"fe",
          1568 => x"0b",
          1569 => x"0c",
          1570 => x"04",
          1571 => x"3f",
          1572 => x"08",
          1573 => x"84",
          1574 => x"04",
          1575 => x"73",
          1576 => x"26",
          1577 => x"10",
          1578 => x"f4",
          1579 => x"08",
          1580 => x"8c",
          1581 => x"3f",
          1582 => x"04",
          1583 => x"51",
          1584 => x"83",
          1585 => x"83",
          1586 => x"ef",
          1587 => x"3d",
          1588 => x"ce",
          1589 => x"9d",
          1590 => x"0d",
          1591 => x"e4",
          1592 => x"3f",
          1593 => x"04",
          1594 => x"51",
          1595 => x"83",
          1596 => x"83",
          1597 => x"ee",
          1598 => x"3d",
          1599 => x"cf",
          1600 => x"f1",
          1601 => x"0d",
          1602 => x"cc",
          1603 => x"3f",
          1604 => x"04",
          1605 => x"51",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ee",
          1609 => x"3d",
          1610 => x"d0",
          1611 => x"c5",
          1612 => x"0d",
          1613 => x"ac",
          1614 => x"3f",
          1615 => x"04",
          1616 => x"51",
          1617 => x"83",
          1618 => x"83",
          1619 => x"ee",
          1620 => x"3d",
          1621 => x"d0",
          1622 => x"99",
          1623 => x"0d",
          1624 => x"f8",
          1625 => x"3f",
          1626 => x"04",
          1627 => x"51",
          1628 => x"83",
          1629 => x"83",
          1630 => x"ed",
          1631 => x"3d",
          1632 => x"d1",
          1633 => x"ed",
          1634 => x"0d",
          1635 => x"b4",
          1636 => x"3f",
          1637 => x"04",
          1638 => x"66",
          1639 => x"80",
          1640 => x"5b",
          1641 => x"79",
          1642 => x"07",
          1643 => x"57",
          1644 => x"57",
          1645 => x"26",
          1646 => x"57",
          1647 => x"70",
          1648 => x"51",
          1649 => x"74",
          1650 => x"81",
          1651 => x"8c",
          1652 => x"58",
          1653 => x"3f",
          1654 => x"08",
          1655 => x"e4",
          1656 => x"80",
          1657 => x"51",
          1658 => x"3f",
          1659 => x"78",
          1660 => x"7b",
          1661 => x"2a",
          1662 => x"57",
          1663 => x"80",
          1664 => x"87",
          1665 => x"08",
          1666 => x"e7",
          1667 => x"38",
          1668 => x"87",
          1669 => x"f5",
          1670 => x"b8",
          1671 => x"83",
          1672 => x"78",
          1673 => x"c0",
          1674 => x"3f",
          1675 => x"e4",
          1676 => x"0d",
          1677 => x"e4",
          1678 => x"98",
          1679 => x"b8",
          1680 => x"96",
          1681 => x"54",
          1682 => x"75",
          1683 => x"82",
          1684 => x"84",
          1685 => x"57",
          1686 => x"08",
          1687 => x"7a",
          1688 => x"2e",
          1689 => x"74",
          1690 => x"57",
          1691 => x"87",
          1692 => x"51",
          1693 => x"84",
          1694 => x"52",
          1695 => x"a7",
          1696 => x"e4",
          1697 => x"d1",
          1698 => x"52",
          1699 => x"51",
          1700 => x"ff",
          1701 => x"3d",
          1702 => x"84",
          1703 => x"33",
          1704 => x"58",
          1705 => x"52",
          1706 => x"ec",
          1707 => x"e4",
          1708 => x"76",
          1709 => x"38",
          1710 => x"8a",
          1711 => x"b8",
          1712 => x"3d",
          1713 => x"04",
          1714 => x"56",
          1715 => x"54",
          1716 => x"53",
          1717 => x"51",
          1718 => x"b8",
          1719 => x"b8",
          1720 => x"3d",
          1721 => x"3d",
          1722 => x"63",
          1723 => x"80",
          1724 => x"73",
          1725 => x"41",
          1726 => x"5f",
          1727 => x"80",
          1728 => x"38",
          1729 => x"d1",
          1730 => x"fe",
          1731 => x"f4",
          1732 => x"3f",
          1733 => x"79",
          1734 => x"7c",
          1735 => x"ed",
          1736 => x"2e",
          1737 => x"73",
          1738 => x"7a",
          1739 => x"38",
          1740 => x"83",
          1741 => x"dd",
          1742 => x"14",
          1743 => x"08",
          1744 => x"51",
          1745 => x"78",
          1746 => x"38",
          1747 => x"51",
          1748 => x"80",
          1749 => x"27",
          1750 => x"75",
          1751 => x"55",
          1752 => x"72",
          1753 => x"38",
          1754 => x"53",
          1755 => x"83",
          1756 => x"74",
          1757 => x"81",
          1758 => x"57",
          1759 => x"88",
          1760 => x"74",
          1761 => x"38",
          1762 => x"08",
          1763 => x"eb",
          1764 => x"16",
          1765 => x"26",
          1766 => x"d2",
          1767 => x"d5",
          1768 => x"79",
          1769 => x"80",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"98",
          1773 => x"76",
          1774 => x"ee",
          1775 => x"2e",
          1776 => x"7b",
          1777 => x"78",
          1778 => x"38",
          1779 => x"b8",
          1780 => x"3d",
          1781 => x"d2",
          1782 => x"ae",
          1783 => x"84",
          1784 => x"53",
          1785 => x"eb",
          1786 => x"74",
          1787 => x"38",
          1788 => x"83",
          1789 => x"dc",
          1790 => x"14",
          1791 => x"08",
          1792 => x"51",
          1793 => x"73",
          1794 => x"c0",
          1795 => x"53",
          1796 => x"df",
          1797 => x"52",
          1798 => x"51",
          1799 => x"82",
          1800 => x"c8",
          1801 => x"a0",
          1802 => x"3f",
          1803 => x"dd",
          1804 => x"39",
          1805 => x"51",
          1806 => x"84",
          1807 => x"c8",
          1808 => x"a0",
          1809 => x"3f",
          1810 => x"fd",
          1811 => x"18",
          1812 => x"27",
          1813 => x"08",
          1814 => x"ec",
          1815 => x"3f",
          1816 => x"d4",
          1817 => x"54",
          1818 => x"84",
          1819 => x"26",
          1820 => x"d8",
          1821 => x"c8",
          1822 => x"51",
          1823 => x"81",
          1824 => x"91",
          1825 => x"d8",
          1826 => x"e4",
          1827 => x"06",
          1828 => x"72",
          1829 => x"ec",
          1830 => x"72",
          1831 => x"09",
          1832 => x"e0",
          1833 => x"fc",
          1834 => x"51",
          1835 => x"84",
          1836 => x"98",
          1837 => x"2c",
          1838 => x"70",
          1839 => x"32",
          1840 => x"72",
          1841 => x"07",
          1842 => x"58",
          1843 => x"53",
          1844 => x"fd",
          1845 => x"51",
          1846 => x"84",
          1847 => x"98",
          1848 => x"2c",
          1849 => x"70",
          1850 => x"32",
          1851 => x"72",
          1852 => x"07",
          1853 => x"58",
          1854 => x"53",
          1855 => x"ff",
          1856 => x"b9",
          1857 => x"84",
          1858 => x"8f",
          1859 => x"fe",
          1860 => x"c0",
          1861 => x"53",
          1862 => x"81",
          1863 => x"3f",
          1864 => x"51",
          1865 => x"80",
          1866 => x"3f",
          1867 => x"70",
          1868 => x"52",
          1869 => x"38",
          1870 => x"70",
          1871 => x"52",
          1872 => x"38",
          1873 => x"70",
          1874 => x"52",
          1875 => x"38",
          1876 => x"70",
          1877 => x"52",
          1878 => x"38",
          1879 => x"70",
          1880 => x"52",
          1881 => x"38",
          1882 => x"70",
          1883 => x"52",
          1884 => x"38",
          1885 => x"70",
          1886 => x"52",
          1887 => x"72",
          1888 => x"06",
          1889 => x"38",
          1890 => x"84",
          1891 => x"81",
          1892 => x"3f",
          1893 => x"51",
          1894 => x"80",
          1895 => x"3f",
          1896 => x"84",
          1897 => x"81",
          1898 => x"3f",
          1899 => x"51",
          1900 => x"80",
          1901 => x"3f",
          1902 => x"81",
          1903 => x"80",
          1904 => x"cb",
          1905 => x"9b",
          1906 => x"d3",
          1907 => x"d4",
          1908 => x"9b",
          1909 => x"87",
          1910 => x"06",
          1911 => x"80",
          1912 => x"38",
          1913 => x"51",
          1914 => x"83",
          1915 => x"9b",
          1916 => x"51",
          1917 => x"72",
          1918 => x"81",
          1919 => x"71",
          1920 => x"f0",
          1921 => x"39",
          1922 => x"80",
          1923 => x"c4",
          1924 => x"3f",
          1925 => x"f4",
          1926 => x"2a",
          1927 => x"51",
          1928 => x"2e",
          1929 => x"ff",
          1930 => x"51",
          1931 => x"83",
          1932 => x"9a",
          1933 => x"51",
          1934 => x"72",
          1935 => x"81",
          1936 => x"71",
          1937 => x"94",
          1938 => x"39",
          1939 => x"bc",
          1940 => x"ec",
          1941 => x"3f",
          1942 => x"b0",
          1943 => x"2a",
          1944 => x"51",
          1945 => x"2e",
          1946 => x"ff",
          1947 => x"51",
          1948 => x"83",
          1949 => x"9a",
          1950 => x"51",
          1951 => x"72",
          1952 => x"81",
          1953 => x"71",
          1954 => x"b8",
          1955 => x"39",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"f0",
          1959 => x"52",
          1960 => x"b5",
          1961 => x"b8",
          1962 => x"ff",
          1963 => x"40",
          1964 => x"2e",
          1965 => x"83",
          1966 => x"e3",
          1967 => x"3d",
          1968 => x"88",
          1969 => x"3f",
          1970 => x"f8",
          1971 => x"7e",
          1972 => x"3f",
          1973 => x"ed",
          1974 => x"81",
          1975 => x"59",
          1976 => x"82",
          1977 => x"81",
          1978 => x"38",
          1979 => x"06",
          1980 => x"2e",
          1981 => x"67",
          1982 => x"79",
          1983 => x"dc",
          1984 => x"5c",
          1985 => x"09",
          1986 => x"38",
          1987 => x"33",
          1988 => x"a0",
          1989 => x"80",
          1990 => x"26",
          1991 => x"90",
          1992 => x"dc",
          1993 => x"52",
          1994 => x"3f",
          1995 => x"08",
          1996 => x"08",
          1997 => x"7b",
          1998 => x"e8",
          1999 => x"b8",
          2000 => x"38",
          2001 => x"5e",
          2002 => x"83",
          2003 => x"1c",
          2004 => x"06",
          2005 => x"7c",
          2006 => x"9a",
          2007 => x"7b",
          2008 => x"dd",
          2009 => x"52",
          2010 => x"92",
          2011 => x"e4",
          2012 => x"b8",
          2013 => x"2e",
          2014 => x"84",
          2015 => x"48",
          2016 => x"80",
          2017 => x"89",
          2018 => x"e4",
          2019 => x"06",
          2020 => x"80",
          2021 => x"38",
          2022 => x"08",
          2023 => x"3f",
          2024 => x"08",
          2025 => x"f3",
          2026 => x"a5",
          2027 => x"7a",
          2028 => x"85",
          2029 => x"24",
          2030 => x"7a",
          2031 => x"e4",
          2032 => x"80",
          2033 => x"8c",
          2034 => x"d5",
          2035 => x"f1",
          2036 => x"b9",
          2037 => x"56",
          2038 => x"54",
          2039 => x"53",
          2040 => x"52",
          2041 => x"ae",
          2042 => x"e4",
          2043 => x"e4",
          2044 => x"30",
          2045 => x"80",
          2046 => x"5b",
          2047 => x"7a",
          2048 => x"38",
          2049 => x"7a",
          2050 => x"80",
          2051 => x"81",
          2052 => x"ff",
          2053 => x"7a",
          2054 => x"7f",
          2055 => x"81",
          2056 => x"7c",
          2057 => x"61",
          2058 => x"e8",
          2059 => x"81",
          2060 => x"83",
          2061 => x"d3",
          2062 => x"48",
          2063 => x"80",
          2064 => x"e8",
          2065 => x"0b",
          2066 => x"33",
          2067 => x"06",
          2068 => x"fd",
          2069 => x"53",
          2070 => x"52",
          2071 => x"51",
          2072 => x"3f",
          2073 => x"08",
          2074 => x"81",
          2075 => x"83",
          2076 => x"84",
          2077 => x"80",
          2078 => x"51",
          2079 => x"3f",
          2080 => x"08",
          2081 => x"38",
          2082 => x"08",
          2083 => x"3f",
          2084 => x"ed",
          2085 => x"81",
          2086 => x"59",
          2087 => x"09",
          2088 => x"d3",
          2089 => x"84",
          2090 => x"82",
          2091 => x"82",
          2092 => x"83",
          2093 => x"83",
          2094 => x"80",
          2095 => x"51",
          2096 => x"67",
          2097 => x"79",
          2098 => x"90",
          2099 => x"63",
          2100 => x"33",
          2101 => x"89",
          2102 => x"38",
          2103 => x"83",
          2104 => x"5a",
          2105 => x"83",
          2106 => x"94",
          2107 => x"e4",
          2108 => x"53",
          2109 => x"ba",
          2110 => x"84",
          2111 => x"b8",
          2112 => x"2e",
          2113 => x"fb",
          2114 => x"70",
          2115 => x"41",
          2116 => x"39",
          2117 => x"51",
          2118 => x"7d",
          2119 => x"e2",
          2120 => x"39",
          2121 => x"56",
          2122 => x"d5",
          2123 => x"53",
          2124 => x"52",
          2125 => x"f2",
          2126 => x"39",
          2127 => x"3f",
          2128 => x"9a",
          2129 => x"f9",
          2130 => x"83",
          2131 => x"3f",
          2132 => x"81",
          2133 => x"fa",
          2134 => x"d5",
          2135 => x"95",
          2136 => x"78",
          2137 => x"d4",
          2138 => x"3f",
          2139 => x"fa",
          2140 => x"3d",
          2141 => x"53",
          2142 => x"51",
          2143 => x"84",
          2144 => x"80",
          2145 => x"38",
          2146 => x"d5",
          2147 => x"fa",
          2148 => x"79",
          2149 => x"e4",
          2150 => x"fa",
          2151 => x"b8",
          2152 => x"83",
          2153 => x"d0",
          2154 => x"95",
          2155 => x"ff",
          2156 => x"ff",
          2157 => x"eb",
          2158 => x"b8",
          2159 => x"2e",
          2160 => x"68",
          2161 => x"a8",
          2162 => x"3f",
          2163 => x"04",
          2164 => x"f4",
          2165 => x"80",
          2166 => x"a8",
          2167 => x"e4",
          2168 => x"f9",
          2169 => x"3d",
          2170 => x"53",
          2171 => x"51",
          2172 => x"84",
          2173 => x"86",
          2174 => x"59",
          2175 => x"78",
          2176 => x"c4",
          2177 => x"3f",
          2178 => x"08",
          2179 => x"52",
          2180 => x"91",
          2181 => x"7e",
          2182 => x"ae",
          2183 => x"38",
          2184 => x"87",
          2185 => x"84",
          2186 => x"59",
          2187 => x"3d",
          2188 => x"53",
          2189 => x"51",
          2190 => x"84",
          2191 => x"80",
          2192 => x"38",
          2193 => x"f0",
          2194 => x"80",
          2195 => x"b4",
          2196 => x"e4",
          2197 => x"38",
          2198 => x"22",
          2199 => x"83",
          2200 => x"cf",
          2201 => x"d4",
          2202 => x"80",
          2203 => x"51",
          2204 => x"7e",
          2205 => x"59",
          2206 => x"f8",
          2207 => x"9f",
          2208 => x"38",
          2209 => x"70",
          2210 => x"39",
          2211 => x"84",
          2212 => x"80",
          2213 => x"f0",
          2214 => x"e4",
          2215 => x"f8",
          2216 => x"3d",
          2217 => x"53",
          2218 => x"51",
          2219 => x"84",
          2220 => x"80",
          2221 => x"38",
          2222 => x"f8",
          2223 => x"80",
          2224 => x"c4",
          2225 => x"e4",
          2226 => x"f7",
          2227 => x"d6",
          2228 => x"b6",
          2229 => x"5d",
          2230 => x"27",
          2231 => x"65",
          2232 => x"33",
          2233 => x"7a",
          2234 => x"38",
          2235 => x"54",
          2236 => x"78",
          2237 => x"f0",
          2238 => x"3f",
          2239 => x"5c",
          2240 => x"1b",
          2241 => x"39",
          2242 => x"84",
          2243 => x"80",
          2244 => x"f4",
          2245 => x"e4",
          2246 => x"f7",
          2247 => x"3d",
          2248 => x"53",
          2249 => x"51",
          2250 => x"84",
          2251 => x"80",
          2252 => x"38",
          2253 => x"f8",
          2254 => x"80",
          2255 => x"c8",
          2256 => x"e4",
          2257 => x"f6",
          2258 => x"d7",
          2259 => x"ba",
          2260 => x"79",
          2261 => x"93",
          2262 => x"79",
          2263 => x"5b",
          2264 => x"65",
          2265 => x"eb",
          2266 => x"ff",
          2267 => x"ff",
          2268 => x"e8",
          2269 => x"b8",
          2270 => x"2e",
          2271 => x"b8",
          2272 => x"11",
          2273 => x"05",
          2274 => x"3f",
          2275 => x"08",
          2276 => x"70",
          2277 => x"83",
          2278 => x"cc",
          2279 => x"d4",
          2280 => x"80",
          2281 => x"51",
          2282 => x"7e",
          2283 => x"59",
          2284 => x"f6",
          2285 => x"9f",
          2286 => x"38",
          2287 => x"49",
          2288 => x"59",
          2289 => x"05",
          2290 => x"68",
          2291 => x"b8",
          2292 => x"11",
          2293 => x"05",
          2294 => x"3f",
          2295 => x"08",
          2296 => x"dd",
          2297 => x"02",
          2298 => x"33",
          2299 => x"81",
          2300 => x"3d",
          2301 => x"53",
          2302 => x"51",
          2303 => x"84",
          2304 => x"ff",
          2305 => x"b9",
          2306 => x"ff",
          2307 => x"ff",
          2308 => x"e6",
          2309 => x"b8",
          2310 => x"2e",
          2311 => x"b8",
          2312 => x"11",
          2313 => x"05",
          2314 => x"3f",
          2315 => x"08",
          2316 => x"8d",
          2317 => x"fe",
          2318 => x"ff",
          2319 => x"e6",
          2320 => x"b8",
          2321 => x"38",
          2322 => x"08",
          2323 => x"a4",
          2324 => x"3f",
          2325 => x"59",
          2326 => x"8f",
          2327 => x"7a",
          2328 => x"05",
          2329 => x"79",
          2330 => x"8a",
          2331 => x"3f",
          2332 => x"b8",
          2333 => x"05",
          2334 => x"3f",
          2335 => x"08",
          2336 => x"80",
          2337 => x"88",
          2338 => x"53",
          2339 => x"08",
          2340 => x"ea",
          2341 => x"b8",
          2342 => x"2e",
          2343 => x"84",
          2344 => x"51",
          2345 => x"f4",
          2346 => x"3d",
          2347 => x"53",
          2348 => x"51",
          2349 => x"84",
          2350 => x"91",
          2351 => x"e8",
          2352 => x"80",
          2353 => x"38",
          2354 => x"08",
          2355 => x"fe",
          2356 => x"ff",
          2357 => x"e5",
          2358 => x"b8",
          2359 => x"38",
          2360 => x"33",
          2361 => x"2e",
          2362 => x"83",
          2363 => x"47",
          2364 => x"f8",
          2365 => x"80",
          2366 => x"8c",
          2367 => x"e4",
          2368 => x"a5",
          2369 => x"5c",
          2370 => x"2e",
          2371 => x"5c",
          2372 => x"70",
          2373 => x"07",
          2374 => x"06",
          2375 => x"79",
          2376 => x"38",
          2377 => x"83",
          2378 => x"83",
          2379 => x"d6",
          2380 => x"55",
          2381 => x"53",
          2382 => x"51",
          2383 => x"83",
          2384 => x"d6",
          2385 => x"f9",
          2386 => x"71",
          2387 => x"84",
          2388 => x"3d",
          2389 => x"53",
          2390 => x"51",
          2391 => x"84",
          2392 => x"80",
          2393 => x"38",
          2394 => x"0c",
          2395 => x"05",
          2396 => x"fe",
          2397 => x"ff",
          2398 => x"e2",
          2399 => x"b8",
          2400 => x"38",
          2401 => x"64",
          2402 => x"ce",
          2403 => x"70",
          2404 => x"23",
          2405 => x"3d",
          2406 => x"53",
          2407 => x"51",
          2408 => x"84",
          2409 => x"80",
          2410 => x"38",
          2411 => x"80",
          2412 => x"7e",
          2413 => x"40",
          2414 => x"b8",
          2415 => x"11",
          2416 => x"05",
          2417 => x"3f",
          2418 => x"08",
          2419 => x"f1",
          2420 => x"3d",
          2421 => x"53",
          2422 => x"51",
          2423 => x"84",
          2424 => x"80",
          2425 => x"38",
          2426 => x"80",
          2427 => x"7c",
          2428 => x"05",
          2429 => x"39",
          2430 => x"f0",
          2431 => x"80",
          2432 => x"80",
          2433 => x"e4",
          2434 => x"81",
          2435 => x"64",
          2436 => x"64",
          2437 => x"46",
          2438 => x"39",
          2439 => x"09",
          2440 => x"9d",
          2441 => x"83",
          2442 => x"80",
          2443 => x"cc",
          2444 => x"c8",
          2445 => x"96",
          2446 => x"7c",
          2447 => x"3f",
          2448 => x"83",
          2449 => x"d4",
          2450 => x"f5",
          2451 => x"fe",
          2452 => x"ff",
          2453 => x"e0",
          2454 => x"b8",
          2455 => x"2e",
          2456 => x"59",
          2457 => x"05",
          2458 => x"82",
          2459 => x"78",
          2460 => x"39",
          2461 => x"33",
          2462 => x"2e",
          2463 => x"83",
          2464 => x"47",
          2465 => x"83",
          2466 => x"5c",
          2467 => x"a1",
          2468 => x"a8",
          2469 => x"b5",
          2470 => x"84",
          2471 => x"3f",
          2472 => x"b6",
          2473 => x"84",
          2474 => x"3f",
          2475 => x"cc",
          2476 => x"ea",
          2477 => x"80",
          2478 => x"83",
          2479 => x"49",
          2480 => x"83",
          2481 => x"d3",
          2482 => x"c6",
          2483 => x"ea",
          2484 => x"80",
          2485 => x"83",
          2486 => x"47",
          2487 => x"83",
          2488 => x"5e",
          2489 => x"9b",
          2490 => x"b8",
          2491 => x"dd",
          2492 => x"eb",
          2493 => x"80",
          2494 => x"83",
          2495 => x"47",
          2496 => x"83",
          2497 => x"5d",
          2498 => x"9b",
          2499 => x"c0",
          2500 => x"b9",
          2501 => x"e6",
          2502 => x"80",
          2503 => x"83",
          2504 => x"47",
          2505 => x"83",
          2506 => x"fc",
          2507 => x"fb",
          2508 => x"f1",
          2509 => x"05",
          2510 => x"39",
          2511 => x"80",
          2512 => x"94",
          2513 => x"94",
          2514 => x"56",
          2515 => x"80",
          2516 => x"da",
          2517 => x"b8",
          2518 => x"2b",
          2519 => x"55",
          2520 => x"52",
          2521 => x"bf",
          2522 => x"b8",
          2523 => x"77",
          2524 => x"94",
          2525 => x"56",
          2526 => x"80",
          2527 => x"da",
          2528 => x"b8",
          2529 => x"2b",
          2530 => x"55",
          2531 => x"52",
          2532 => x"93",
          2533 => x"b8",
          2534 => x"77",
          2535 => x"83",
          2536 => x"94",
          2537 => x"80",
          2538 => x"c0",
          2539 => x"81",
          2540 => x"81",
          2541 => x"83",
          2542 => x"a1",
          2543 => x"5e",
          2544 => x"0b",
          2545 => x"88",
          2546 => x"72",
          2547 => x"c8",
          2548 => x"f4",
          2549 => x"3f",
          2550 => x"ba",
          2551 => x"fc",
          2552 => x"a0",
          2553 => x"a4",
          2554 => x"3f",
          2555 => x"70",
          2556 => x"94",
          2557 => x"d2",
          2558 => x"d2",
          2559 => x"15",
          2560 => x"d2",
          2561 => x"82",
          2562 => x"3f",
          2563 => x"80",
          2564 => x"0d",
          2565 => x"56",
          2566 => x"52",
          2567 => x"2e",
          2568 => x"74",
          2569 => x"ff",
          2570 => x"70",
          2571 => x"81",
          2572 => x"81",
          2573 => x"70",
          2574 => x"53",
          2575 => x"a0",
          2576 => x"71",
          2577 => x"54",
          2578 => x"81",
          2579 => x"52",
          2580 => x"80",
          2581 => x"72",
          2582 => x"ff",
          2583 => x"54",
          2584 => x"83",
          2585 => x"70",
          2586 => x"38",
          2587 => x"86",
          2588 => x"52",
          2589 => x"73",
          2590 => x"52",
          2591 => x"2e",
          2592 => x"83",
          2593 => x"70",
          2594 => x"30",
          2595 => x"76",
          2596 => x"53",
          2597 => x"88",
          2598 => x"70",
          2599 => x"34",
          2600 => x"74",
          2601 => x"b8",
          2602 => x"3d",
          2603 => x"80",
          2604 => x"73",
          2605 => x"be",
          2606 => x"52",
          2607 => x"70",
          2608 => x"53",
          2609 => x"a2",
          2610 => x"81",
          2611 => x"81",
          2612 => x"75",
          2613 => x"81",
          2614 => x"06",
          2615 => x"dc",
          2616 => x"0d",
          2617 => x"08",
          2618 => x"0b",
          2619 => x"0c",
          2620 => x"04",
          2621 => x"05",
          2622 => x"db",
          2623 => x"b8",
          2624 => x"2e",
          2625 => x"84",
          2626 => x"86",
          2627 => x"fc",
          2628 => x"82",
          2629 => x"05",
          2630 => x"52",
          2631 => x"81",
          2632 => x"13",
          2633 => x"54",
          2634 => x"9e",
          2635 => x"38",
          2636 => x"51",
          2637 => x"97",
          2638 => x"38",
          2639 => x"54",
          2640 => x"bb",
          2641 => x"38",
          2642 => x"55",
          2643 => x"bb",
          2644 => x"38",
          2645 => x"55",
          2646 => x"87",
          2647 => x"d9",
          2648 => x"22",
          2649 => x"73",
          2650 => x"80",
          2651 => x"0b",
          2652 => x"9c",
          2653 => x"87",
          2654 => x"0c",
          2655 => x"87",
          2656 => x"0c",
          2657 => x"87",
          2658 => x"0c",
          2659 => x"87",
          2660 => x"0c",
          2661 => x"87",
          2662 => x"0c",
          2663 => x"87",
          2664 => x"0c",
          2665 => x"98",
          2666 => x"87",
          2667 => x"0c",
          2668 => x"c0",
          2669 => x"80",
          2670 => x"b8",
          2671 => x"3d",
          2672 => x"3d",
          2673 => x"87",
          2674 => x"5d",
          2675 => x"87",
          2676 => x"08",
          2677 => x"23",
          2678 => x"b8",
          2679 => x"82",
          2680 => x"c0",
          2681 => x"5a",
          2682 => x"34",
          2683 => x"b0",
          2684 => x"84",
          2685 => x"c0",
          2686 => x"5a",
          2687 => x"34",
          2688 => x"a8",
          2689 => x"86",
          2690 => x"c0",
          2691 => x"5c",
          2692 => x"23",
          2693 => x"a0",
          2694 => x"8a",
          2695 => x"7d",
          2696 => x"ff",
          2697 => x"7b",
          2698 => x"06",
          2699 => x"33",
          2700 => x"33",
          2701 => x"33",
          2702 => x"33",
          2703 => x"33",
          2704 => x"ff",
          2705 => x"83",
          2706 => x"ff",
          2707 => x"8f",
          2708 => x"fe",
          2709 => x"93",
          2710 => x"72",
          2711 => x"38",
          2712 => x"e8",
          2713 => x"b8",
          2714 => x"2b",
          2715 => x"51",
          2716 => x"2e",
          2717 => x"86",
          2718 => x"2e",
          2719 => x"84",
          2720 => x"84",
          2721 => x"72",
          2722 => x"89",
          2723 => x"e4",
          2724 => x"70",
          2725 => x"52",
          2726 => x"09",
          2727 => x"38",
          2728 => x"e7",
          2729 => x"b8",
          2730 => x"2b",
          2731 => x"51",
          2732 => x"2e",
          2733 => x"39",
          2734 => x"80",
          2735 => x"71",
          2736 => x"81",
          2737 => x"cd",
          2738 => x"e4",
          2739 => x"70",
          2740 => x"52",
          2741 => x"eb",
          2742 => x"07",
          2743 => x"52",
          2744 => x"db",
          2745 => x"b8",
          2746 => x"3d",
          2747 => x"3d",
          2748 => x"05",
          2749 => x"9c",
          2750 => x"ff",
          2751 => x"55",
          2752 => x"80",
          2753 => x"c0",
          2754 => x"70",
          2755 => x"81",
          2756 => x"52",
          2757 => x"8c",
          2758 => x"2a",
          2759 => x"51",
          2760 => x"38",
          2761 => x"81",
          2762 => x"80",
          2763 => x"71",
          2764 => x"06",
          2765 => x"38",
          2766 => x"06",
          2767 => x"94",
          2768 => x"80",
          2769 => x"87",
          2770 => x"52",
          2771 => x"74",
          2772 => x"0c",
          2773 => x"04",
          2774 => x"70",
          2775 => x"51",
          2776 => x"72",
          2777 => x"06",
          2778 => x"2e",
          2779 => x"93",
          2780 => x"52",
          2781 => x"c0",
          2782 => x"94",
          2783 => x"96",
          2784 => x"06",
          2785 => x"70",
          2786 => x"39",
          2787 => x"02",
          2788 => x"70",
          2789 => x"2a",
          2790 => x"70",
          2791 => x"34",
          2792 => x"04",
          2793 => x"78",
          2794 => x"33",
          2795 => x"57",
          2796 => x"80",
          2797 => x"15",
          2798 => x"33",
          2799 => x"06",
          2800 => x"71",
          2801 => x"ff",
          2802 => x"94",
          2803 => x"96",
          2804 => x"06",
          2805 => x"70",
          2806 => x"38",
          2807 => x"70",
          2808 => x"51",
          2809 => x"72",
          2810 => x"06",
          2811 => x"2e",
          2812 => x"93",
          2813 => x"52",
          2814 => x"75",
          2815 => x"51",
          2816 => x"80",
          2817 => x"2e",
          2818 => x"c0",
          2819 => x"73",
          2820 => x"17",
          2821 => x"57",
          2822 => x"38",
          2823 => x"e4",
          2824 => x"0d",
          2825 => x"2a",
          2826 => x"51",
          2827 => x"38",
          2828 => x"81",
          2829 => x"80",
          2830 => x"71",
          2831 => x"06",
          2832 => x"2e",
          2833 => x"87",
          2834 => x"08",
          2835 => x"70",
          2836 => x"54",
          2837 => x"38",
          2838 => x"3d",
          2839 => x"9e",
          2840 => x"9c",
          2841 => x"52",
          2842 => x"2e",
          2843 => x"87",
          2844 => x"08",
          2845 => x"0c",
          2846 => x"a8",
          2847 => x"a4",
          2848 => x"9e",
          2849 => x"f1",
          2850 => x"c0",
          2851 => x"83",
          2852 => x"87",
          2853 => x"08",
          2854 => x"0c",
          2855 => x"a0",
          2856 => x"b4",
          2857 => x"9e",
          2858 => x"f1",
          2859 => x"c0",
          2860 => x"83",
          2861 => x"87",
          2862 => x"08",
          2863 => x"0c",
          2864 => x"b8",
          2865 => x"c4",
          2866 => x"9e",
          2867 => x"f1",
          2868 => x"c0",
          2869 => x"83",
          2870 => x"87",
          2871 => x"08",
          2872 => x"0c",
          2873 => x"80",
          2874 => x"83",
          2875 => x"87",
          2876 => x"08",
          2877 => x"0c",
          2878 => x"88",
          2879 => x"dc",
          2880 => x"9e",
          2881 => x"f1",
          2882 => x"0b",
          2883 => x"34",
          2884 => x"c0",
          2885 => x"70",
          2886 => x"06",
          2887 => x"70",
          2888 => x"71",
          2889 => x"34",
          2890 => x"c0",
          2891 => x"70",
          2892 => x"06",
          2893 => x"70",
          2894 => x"38",
          2895 => x"83",
          2896 => x"80",
          2897 => x"9e",
          2898 => x"90",
          2899 => x"51",
          2900 => x"80",
          2901 => x"81",
          2902 => x"f1",
          2903 => x"0b",
          2904 => x"90",
          2905 => x"80",
          2906 => x"52",
          2907 => x"2e",
          2908 => x"52",
          2909 => x"e8",
          2910 => x"87",
          2911 => x"08",
          2912 => x"80",
          2913 => x"52",
          2914 => x"83",
          2915 => x"71",
          2916 => x"34",
          2917 => x"c0",
          2918 => x"70",
          2919 => x"06",
          2920 => x"70",
          2921 => x"38",
          2922 => x"83",
          2923 => x"80",
          2924 => x"9e",
          2925 => x"84",
          2926 => x"51",
          2927 => x"80",
          2928 => x"81",
          2929 => x"f1",
          2930 => x"0b",
          2931 => x"90",
          2932 => x"80",
          2933 => x"52",
          2934 => x"2e",
          2935 => x"52",
          2936 => x"ec",
          2937 => x"87",
          2938 => x"08",
          2939 => x"80",
          2940 => x"52",
          2941 => x"83",
          2942 => x"71",
          2943 => x"34",
          2944 => x"c0",
          2945 => x"70",
          2946 => x"06",
          2947 => x"70",
          2948 => x"38",
          2949 => x"83",
          2950 => x"80",
          2951 => x"9e",
          2952 => x"a0",
          2953 => x"52",
          2954 => x"2e",
          2955 => x"52",
          2956 => x"ef",
          2957 => x"9e",
          2958 => x"80",
          2959 => x"2a",
          2960 => x"83",
          2961 => x"80",
          2962 => x"9e",
          2963 => x"84",
          2964 => x"52",
          2965 => x"2e",
          2966 => x"52",
          2967 => x"f1",
          2968 => x"9e",
          2969 => x"f0",
          2970 => x"2a",
          2971 => x"83",
          2972 => x"80",
          2973 => x"9e",
          2974 => x"88",
          2975 => x"52",
          2976 => x"83",
          2977 => x"71",
          2978 => x"34",
          2979 => x"90",
          2980 => x"51",
          2981 => x"f4",
          2982 => x"0d",
          2983 => x"fd",
          2984 => x"3d",
          2985 => x"a0",
          2986 => x"de",
          2987 => x"e4",
          2988 => x"86",
          2989 => x"d8",
          2990 => x"b9",
          2991 => x"e6",
          2992 => x"85",
          2993 => x"f1",
          2994 => x"73",
          2995 => x"83",
          2996 => x"56",
          2997 => x"38",
          2998 => x"33",
          2999 => x"ff",
          3000 => x"ea",
          3001 => x"84",
          3002 => x"f1",
          3003 => x"75",
          3004 => x"83",
          3005 => x"54",
          3006 => x"38",
          3007 => x"33",
          3008 => x"ed",
          3009 => x"e5",
          3010 => x"83",
          3011 => x"f1",
          3012 => x"73",
          3013 => x"83",
          3014 => x"55",
          3015 => x"38",
          3016 => x"33",
          3017 => x"f4",
          3018 => x"ee",
          3019 => x"81",
          3020 => x"d8",
          3021 => x"bd",
          3022 => x"c8",
          3023 => x"d8",
          3024 => x"b5",
          3025 => x"f1",
          3026 => x"83",
          3027 => x"ff",
          3028 => x"83",
          3029 => x"52",
          3030 => x"51",
          3031 => x"3f",
          3032 => x"51",
          3033 => x"83",
          3034 => x"52",
          3035 => x"51",
          3036 => x"3f",
          3037 => x"08",
          3038 => x"c0",
          3039 => x"ca",
          3040 => x"b8",
          3041 => x"84",
          3042 => x"71",
          3043 => x"84",
          3044 => x"52",
          3045 => x"51",
          3046 => x"3f",
          3047 => x"33",
          3048 => x"c3",
          3049 => x"e6",
          3050 => x"8a",
          3051 => x"c3",
          3052 => x"3d",
          3053 => x"f1",
          3054 => x"bd",
          3055 => x"75",
          3056 => x"3f",
          3057 => x"08",
          3058 => x"29",
          3059 => x"54",
          3060 => x"e4",
          3061 => x"da",
          3062 => x"b4",
          3063 => x"51",
          3064 => x"87",
          3065 => x"83",
          3066 => x"56",
          3067 => x"52",
          3068 => x"b3",
          3069 => x"e4",
          3070 => x"c0",
          3071 => x"31",
          3072 => x"b8",
          3073 => x"83",
          3074 => x"ff",
          3075 => x"83",
          3076 => x"55",
          3077 => x"ff",
          3078 => x"9a",
          3079 => x"84",
          3080 => x"3f",
          3081 => x"51",
          3082 => x"83",
          3083 => x"52",
          3084 => x"51",
          3085 => x"3f",
          3086 => x"08",
          3087 => x"80",
          3088 => x"c6",
          3089 => x"d0",
          3090 => x"d9",
          3091 => x"b3",
          3092 => x"d9",
          3093 => x"9d",
          3094 => x"d4",
          3095 => x"d9",
          3096 => x"b3",
          3097 => x"f1",
          3098 => x"bd",
          3099 => x"75",
          3100 => x"3f",
          3101 => x"08",
          3102 => x"29",
          3103 => x"54",
          3104 => x"e4",
          3105 => x"da",
          3106 => x"b2",
          3107 => x"f1",
          3108 => x"74",
          3109 => x"8d",
          3110 => x"39",
          3111 => x"51",
          3112 => x"3f",
          3113 => x"33",
          3114 => x"2e",
          3115 => x"fe",
          3116 => x"db",
          3117 => x"bf",
          3118 => x"f1",
          3119 => x"75",
          3120 => x"e5",
          3121 => x"83",
          3122 => x"ff",
          3123 => x"83",
          3124 => x"55",
          3125 => x"fc",
          3126 => x"39",
          3127 => x"51",
          3128 => x"3f",
          3129 => x"33",
          3130 => x"2e",
          3131 => x"d7",
          3132 => x"f2",
          3133 => x"db",
          3134 => x"b2",
          3135 => x"f1",
          3136 => x"75",
          3137 => x"86",
          3138 => x"83",
          3139 => x"52",
          3140 => x"51",
          3141 => x"3f",
          3142 => x"33",
          3143 => x"2e",
          3144 => x"cd",
          3145 => x"f0",
          3146 => x"dc",
          3147 => x"b1",
          3148 => x"f1",
          3149 => x"73",
          3150 => x"c0",
          3151 => x"83",
          3152 => x"83",
          3153 => x"11",
          3154 => x"dc",
          3155 => x"b1",
          3156 => x"f1",
          3157 => x"75",
          3158 => x"97",
          3159 => x"83",
          3160 => x"83",
          3161 => x"11",
          3162 => x"dc",
          3163 => x"b1",
          3164 => x"f1",
          3165 => x"73",
          3166 => x"ee",
          3167 => x"83",
          3168 => x"83",
          3169 => x"11",
          3170 => x"dc",
          3171 => x"b0",
          3172 => x"f1",
          3173 => x"74",
          3174 => x"c5",
          3175 => x"83",
          3176 => x"83",
          3177 => x"11",
          3178 => x"dc",
          3179 => x"b0",
          3180 => x"f1",
          3181 => x"75",
          3182 => x"9c",
          3183 => x"83",
          3184 => x"83",
          3185 => x"11",
          3186 => x"dd",
          3187 => x"b0",
          3188 => x"f1",
          3189 => x"73",
          3190 => x"f3",
          3191 => x"83",
          3192 => x"ff",
          3193 => x"83",
          3194 => x"ff",
          3195 => x"83",
          3196 => x"55",
          3197 => x"f9",
          3198 => x"39",
          3199 => x"02",
          3200 => x"52",
          3201 => x"8c",
          3202 => x"10",
          3203 => x"05",
          3204 => x"04",
          3205 => x"51",
          3206 => x"3f",
          3207 => x"04",
          3208 => x"51",
          3209 => x"3f",
          3210 => x"04",
          3211 => x"51",
          3212 => x"3f",
          3213 => x"04",
          3214 => x"51",
          3215 => x"3f",
          3216 => x"04",
          3217 => x"51",
          3218 => x"3f",
          3219 => x"04",
          3220 => x"51",
          3221 => x"3f",
          3222 => x"04",
          3223 => x"0c",
          3224 => x"87",
          3225 => x"0c",
          3226 => x"f8",
          3227 => x"96",
          3228 => x"d9",
          3229 => x"3d",
          3230 => x"08",
          3231 => x"70",
          3232 => x"52",
          3233 => x"08",
          3234 => x"82",
          3235 => x"e4",
          3236 => x"38",
          3237 => x"ff",
          3238 => x"d0",
          3239 => x"80",
          3240 => x"51",
          3241 => x"3f",
          3242 => x"08",
          3243 => x"38",
          3244 => x"f6",
          3245 => x"e4",
          3246 => x"57",
          3247 => x"84",
          3248 => x"25",
          3249 => x"b8",
          3250 => x"05",
          3251 => x"55",
          3252 => x"74",
          3253 => x"70",
          3254 => x"2a",
          3255 => x"78",
          3256 => x"38",
          3257 => x"38",
          3258 => x"08",
          3259 => x"53",
          3260 => x"9a",
          3261 => x"e4",
          3262 => x"78",
          3263 => x"38",
          3264 => x"e4",
          3265 => x"0d",
          3266 => x"98",
          3267 => x"fa",
          3268 => x"2e",
          3269 => x"e8",
          3270 => x"79",
          3271 => x"3f",
          3272 => x"86",
          3273 => x"08",
          3274 => x"e4",
          3275 => x"76",
          3276 => x"c4",
          3277 => x"d2",
          3278 => x"84",
          3279 => x"a9",
          3280 => x"d8",
          3281 => x"3d",
          3282 => x"08",
          3283 => x"72",
          3284 => x"5a",
          3285 => x"2e",
          3286 => x"80",
          3287 => x"59",
          3288 => x"10",
          3289 => x"d8",
          3290 => x"52",
          3291 => x"ba",
          3292 => x"e4",
          3293 => x"52",
          3294 => x"c0",
          3295 => x"b8",
          3296 => x"38",
          3297 => x"54",
          3298 => x"81",
          3299 => x"82",
          3300 => x"81",
          3301 => x"ff",
          3302 => x"82",
          3303 => x"38",
          3304 => x"84",
          3305 => x"aa",
          3306 => x"81",
          3307 => x"3d",
          3308 => x"53",
          3309 => x"51",
          3310 => x"84",
          3311 => x"80",
          3312 => x"ff",
          3313 => x"52",
          3314 => x"a7",
          3315 => x"e4",
          3316 => x"06",
          3317 => x"2e",
          3318 => x"16",
          3319 => x"06",
          3320 => x"76",
          3321 => x"38",
          3322 => x"78",
          3323 => x"56",
          3324 => x"fe",
          3325 => x"15",
          3326 => x"33",
          3327 => x"a0",
          3328 => x"06",
          3329 => x"75",
          3330 => x"38",
          3331 => x"3d",
          3332 => x"cd",
          3333 => x"b8",
          3334 => x"83",
          3335 => x"52",
          3336 => x"ea",
          3337 => x"e4",
          3338 => x"38",
          3339 => x"08",
          3340 => x"52",
          3341 => x"ce",
          3342 => x"b8",
          3343 => x"2e",
          3344 => x"51",
          3345 => x"3f",
          3346 => x"08",
          3347 => x"84",
          3348 => x"25",
          3349 => x"b8",
          3350 => x"05",
          3351 => x"55",
          3352 => x"77",
          3353 => x"81",
          3354 => x"8c",
          3355 => x"ab",
          3356 => x"ff",
          3357 => x"06",
          3358 => x"81",
          3359 => x"e4",
          3360 => x"0d",
          3361 => x"0d",
          3362 => x"b7",
          3363 => x"3d",
          3364 => x"5c",
          3365 => x"3d",
          3366 => x"d4",
          3367 => x"d0",
          3368 => x"74",
          3369 => x"83",
          3370 => x"56",
          3371 => x"2e",
          3372 => x"77",
          3373 => x"8d",
          3374 => x"77",
          3375 => x"78",
          3376 => x"77",
          3377 => x"fd",
          3378 => x"b4",
          3379 => x"80",
          3380 => x"3f",
          3381 => x"08",
          3382 => x"98",
          3383 => x"79",
          3384 => x"38",
          3385 => x"06",
          3386 => x"33",
          3387 => x"70",
          3388 => x"d0",
          3389 => x"98",
          3390 => x"2c",
          3391 => x"05",
          3392 => x"83",
          3393 => x"70",
          3394 => x"33",
          3395 => x"5d",
          3396 => x"58",
          3397 => x"57",
          3398 => x"80",
          3399 => x"75",
          3400 => x"38",
          3401 => x"0a",
          3402 => x"0a",
          3403 => x"2c",
          3404 => x"76",
          3405 => x"38",
          3406 => x"70",
          3407 => x"57",
          3408 => x"dd",
          3409 => x"42",
          3410 => x"25",
          3411 => x"dd",
          3412 => x"18",
          3413 => x"41",
          3414 => x"81",
          3415 => x"80",
          3416 => x"75",
          3417 => x"34",
          3418 => x"80",
          3419 => x"38",
          3420 => x"98",
          3421 => x"2c",
          3422 => x"33",
          3423 => x"70",
          3424 => x"98",
          3425 => x"82",
          3426 => x"f0",
          3427 => x"53",
          3428 => x"5d",
          3429 => x"78",
          3430 => x"38",
          3431 => x"a0",
          3432 => x"39",
          3433 => x"ff",
          3434 => x"81",
          3435 => x"81",
          3436 => x"70",
          3437 => x"81",
          3438 => x"57",
          3439 => x"26",
          3440 => x"75",
          3441 => x"82",
          3442 => x"80",
          3443 => x"f0",
          3444 => x"57",
          3445 => x"ce",
          3446 => x"ec",
          3447 => x"70",
          3448 => x"78",
          3449 => x"bc",
          3450 => x"2e",
          3451 => x"fe",
          3452 => x"57",
          3453 => x"fe",
          3454 => x"e7",
          3455 => x"fd",
          3456 => x"57",
          3457 => x"38",
          3458 => x"a0",
          3459 => x"d0",
          3460 => x"7e",
          3461 => x"0c",
          3462 => x"95",
          3463 => x"38",
          3464 => x"83",
          3465 => x"57",
          3466 => x"83",
          3467 => x"08",
          3468 => x"0b",
          3469 => x"34",
          3470 => x"d0",
          3471 => x"39",
          3472 => x"33",
          3473 => x"2e",
          3474 => x"84",
          3475 => x"52",
          3476 => x"b6",
          3477 => x"d0",
          3478 => x"05",
          3479 => x"d0",
          3480 => x"eb",
          3481 => x"a8",
          3482 => x"ff",
          3483 => x"a4",
          3484 => x"55",
          3485 => x"fc",
          3486 => x"d4",
          3487 => x"81",
          3488 => x"84",
          3489 => x"7b",
          3490 => x"52",
          3491 => x"e0",
          3492 => x"39",
          3493 => x"8b",
          3494 => x"10",
          3495 => x"80",
          3496 => x"57",
          3497 => x"83",
          3498 => x"d0",
          3499 => x"7c",
          3500 => x"a4",
          3501 => x"a8",
          3502 => x"74",
          3503 => x"38",
          3504 => x"08",
          3505 => x"ff",
          3506 => x"84",
          3507 => x"52",
          3508 => x"b5",
          3509 => x"d4",
          3510 => x"88",
          3511 => x"90",
          3512 => x"a8",
          3513 => x"5b",
          3514 => x"a8",
          3515 => x"ff",
          3516 => x"cc",
          3517 => x"ff",
          3518 => x"75",
          3519 => x"34",
          3520 => x"7c",
          3521 => x"f2",
          3522 => x"75",
          3523 => x"7c",
          3524 => x"f1",
          3525 => x"11",
          3526 => x"75",
          3527 => x"74",
          3528 => x"80",
          3529 => x"38",
          3530 => x"b7",
          3531 => x"b8",
          3532 => x"d0",
          3533 => x"b8",
          3534 => x"ff",
          3535 => x"53",
          3536 => x"51",
          3537 => x"3f",
          3538 => x"33",
          3539 => x"33",
          3540 => x"80",
          3541 => x"38",
          3542 => x"08",
          3543 => x"ff",
          3544 => x"84",
          3545 => x"52",
          3546 => x"b4",
          3547 => x"d4",
          3548 => x"88",
          3549 => x"f8",
          3550 => x"a8",
          3551 => x"55",
          3552 => x"a8",
          3553 => x"ff",
          3554 => x"39",
          3555 => x"33",
          3556 => x"06",
          3557 => x"33",
          3558 => x"75",
          3559 => x"af",
          3560 => x"c8",
          3561 => x"15",
          3562 => x"d0",
          3563 => x"16",
          3564 => x"55",
          3565 => x"3f",
          3566 => x"33",
          3567 => x"06",
          3568 => x"33",
          3569 => x"75",
          3570 => x"83",
          3571 => x"c8",
          3572 => x"15",
          3573 => x"d0",
          3574 => x"16",
          3575 => x"55",
          3576 => x"3f",
          3577 => x"33",
          3578 => x"06",
          3579 => x"33",
          3580 => x"77",
          3581 => x"a9",
          3582 => x"39",
          3583 => x"33",
          3584 => x"33",
          3585 => x"76",
          3586 => x"38",
          3587 => x"7a",
          3588 => x"34",
          3589 => x"70",
          3590 => x"81",
          3591 => x"57",
          3592 => x"24",
          3593 => x"84",
          3594 => x"52",
          3595 => x"b2",
          3596 => x"d0",
          3597 => x"98",
          3598 => x"2c",
          3599 => x"33",
          3600 => x"41",
          3601 => x"f9",
          3602 => x"d4",
          3603 => x"88",
          3604 => x"9c",
          3605 => x"80",
          3606 => x"80",
          3607 => x"98",
          3608 => x"a4",
          3609 => x"5a",
          3610 => x"f8",
          3611 => x"d4",
          3612 => x"88",
          3613 => x"f8",
          3614 => x"80",
          3615 => x"80",
          3616 => x"98",
          3617 => x"a4",
          3618 => x"5a",
          3619 => x"ff",
          3620 => x"bb",
          3621 => x"58",
          3622 => x"78",
          3623 => x"c8",
          3624 => x"33",
          3625 => x"c8",
          3626 => x"80",
          3627 => x"80",
          3628 => x"98",
          3629 => x"a4",
          3630 => x"55",
          3631 => x"fe",
          3632 => x"16",
          3633 => x"33",
          3634 => x"d4",
          3635 => x"77",
          3636 => x"b1",
          3637 => x"81",
          3638 => x"81",
          3639 => x"70",
          3640 => x"d0",
          3641 => x"57",
          3642 => x"24",
          3643 => x"fe",
          3644 => x"d0",
          3645 => x"74",
          3646 => x"d3",
          3647 => x"c8",
          3648 => x"51",
          3649 => x"3f",
          3650 => x"33",
          3651 => x"76",
          3652 => x"34",
          3653 => x"06",
          3654 => x"84",
          3655 => x"7c",
          3656 => x"7f",
          3657 => x"c8",
          3658 => x"51",
          3659 => x"3f",
          3660 => x"52",
          3661 => x"8b",
          3662 => x"e4",
          3663 => x"06",
          3664 => x"cf",
          3665 => x"a4",
          3666 => x"80",
          3667 => x"38",
          3668 => x"33",
          3669 => x"83",
          3670 => x"70",
          3671 => x"56",
          3672 => x"38",
          3673 => x"87",
          3674 => x"f1",
          3675 => x"18",
          3676 => x"5b",
          3677 => x"3f",
          3678 => x"08",
          3679 => x"f2",
          3680 => x"10",
          3681 => x"fc",
          3682 => x"57",
          3683 => x"8b",
          3684 => x"f2",
          3685 => x"75",
          3686 => x"38",
          3687 => x"33",
          3688 => x"2e",
          3689 => x"80",
          3690 => x"a8",
          3691 => x"84",
          3692 => x"7b",
          3693 => x"0c",
          3694 => x"04",
          3695 => x"33",
          3696 => x"2e",
          3697 => x"d4",
          3698 => x"88",
          3699 => x"a0",
          3700 => x"c8",
          3701 => x"51",
          3702 => x"3f",
          3703 => x"08",
          3704 => x"ff",
          3705 => x"84",
          3706 => x"ff",
          3707 => x"84",
          3708 => x"75",
          3709 => x"55",
          3710 => x"83",
          3711 => x"ff",
          3712 => x"80",
          3713 => x"a8",
          3714 => x"84",
          3715 => x"f5",
          3716 => x"7c",
          3717 => x"81",
          3718 => x"d0",
          3719 => x"74",
          3720 => x"38",
          3721 => x"08",
          3722 => x"ff",
          3723 => x"84",
          3724 => x"52",
          3725 => x"ae",
          3726 => x"d4",
          3727 => x"88",
          3728 => x"ac",
          3729 => x"a8",
          3730 => x"5d",
          3731 => x"a8",
          3732 => x"ff",
          3733 => x"cc",
          3734 => x"e0",
          3735 => x"aa",
          3736 => x"84",
          3737 => x"80",
          3738 => x"a4",
          3739 => x"b8",
          3740 => x"3d",
          3741 => x"d0",
          3742 => x"81",
          3743 => x"56",
          3744 => x"f4",
          3745 => x"d0",
          3746 => x"05",
          3747 => x"d0",
          3748 => x"16",
          3749 => x"d0",
          3750 => x"d4",
          3751 => x"88",
          3752 => x"cc",
          3753 => x"a8",
          3754 => x"2b",
          3755 => x"84",
          3756 => x"5a",
          3757 => x"76",
          3758 => x"ef",
          3759 => x"c8",
          3760 => x"51",
          3761 => x"3f",
          3762 => x"33",
          3763 => x"70",
          3764 => x"d0",
          3765 => x"57",
          3766 => x"7a",
          3767 => x"38",
          3768 => x"08",
          3769 => x"ff",
          3770 => x"74",
          3771 => x"29",
          3772 => x"05",
          3773 => x"84",
          3774 => x"5b",
          3775 => x"79",
          3776 => x"38",
          3777 => x"08",
          3778 => x"ff",
          3779 => x"74",
          3780 => x"29",
          3781 => x"05",
          3782 => x"84",
          3783 => x"5b",
          3784 => x"75",
          3785 => x"38",
          3786 => x"7b",
          3787 => x"17",
          3788 => x"84",
          3789 => x"52",
          3790 => x"ff",
          3791 => x"75",
          3792 => x"29",
          3793 => x"05",
          3794 => x"84",
          3795 => x"43",
          3796 => x"61",
          3797 => x"38",
          3798 => x"81",
          3799 => x"34",
          3800 => x"08",
          3801 => x"51",
          3802 => x"3f",
          3803 => x"0a",
          3804 => x"0a",
          3805 => x"2c",
          3806 => x"33",
          3807 => x"60",
          3808 => x"a7",
          3809 => x"39",
          3810 => x"33",
          3811 => x"06",
          3812 => x"60",
          3813 => x"38",
          3814 => x"33",
          3815 => x"27",
          3816 => x"98",
          3817 => x"2c",
          3818 => x"76",
          3819 => x"7b",
          3820 => x"33",
          3821 => x"75",
          3822 => x"29",
          3823 => x"05",
          3824 => x"84",
          3825 => x"52",
          3826 => x"78",
          3827 => x"81",
          3828 => x"84",
          3829 => x"77",
          3830 => x"7c",
          3831 => x"3d",
          3832 => x"84",
          3833 => x"57",
          3834 => x"8b",
          3835 => x"56",
          3836 => x"a4",
          3837 => x"84",
          3838 => x"70",
          3839 => x"29",
          3840 => x"05",
          3841 => x"79",
          3842 => x"44",
          3843 => x"60",
          3844 => x"ef",
          3845 => x"2b",
          3846 => x"78",
          3847 => x"5c",
          3848 => x"7a",
          3849 => x"38",
          3850 => x"08",
          3851 => x"ff",
          3852 => x"75",
          3853 => x"29",
          3854 => x"05",
          3855 => x"84",
          3856 => x"57",
          3857 => x"75",
          3858 => x"38",
          3859 => x"08",
          3860 => x"ff",
          3861 => x"75",
          3862 => x"29",
          3863 => x"05",
          3864 => x"84",
          3865 => x"57",
          3866 => x"76",
          3867 => x"38",
          3868 => x"83",
          3869 => x"56",
          3870 => x"f4",
          3871 => x"51",
          3872 => x"3f",
          3873 => x"08",
          3874 => x"34",
          3875 => x"08",
          3876 => x"81",
          3877 => x"52",
          3878 => x"ad",
          3879 => x"d0",
          3880 => x"d0",
          3881 => x"56",
          3882 => x"f4",
          3883 => x"d4",
          3884 => x"88",
          3885 => x"b8",
          3886 => x"c8",
          3887 => x"51",
          3888 => x"3f",
          3889 => x"08",
          3890 => x"ff",
          3891 => x"84",
          3892 => x"ff",
          3893 => x"84",
          3894 => x"7a",
          3895 => x"55",
          3896 => x"51",
          3897 => x"3f",
          3898 => x"08",
          3899 => x"0c",
          3900 => x"08",
          3901 => x"76",
          3902 => x"34",
          3903 => x"38",
          3904 => x"84",
          3905 => x"52",
          3906 => x"33",
          3907 => x"a8",
          3908 => x"81",
          3909 => x"81",
          3910 => x"70",
          3911 => x"d0",
          3912 => x"57",
          3913 => x"24",
          3914 => x"d0",
          3915 => x"98",
          3916 => x"2c",
          3917 => x"06",
          3918 => x"58",
          3919 => x"ef",
          3920 => x"e4",
          3921 => x"d0",
          3922 => x"ee",
          3923 => x"f1",
          3924 => x"56",
          3925 => x"74",
          3926 => x"16",
          3927 => x"56",
          3928 => x"f0",
          3929 => x"83",
          3930 => x"83",
          3931 => x"55",
          3932 => x"ee",
          3933 => x"51",
          3934 => x"3f",
          3935 => x"08",
          3936 => x"fe",
          3937 => x"83",
          3938 => x"93",
          3939 => x"5f",
          3940 => x"39",
          3941 => x"d9",
          3942 => x"77",
          3943 => x"84",
          3944 => x"75",
          3945 => x"ac",
          3946 => x"39",
          3947 => x"aa",
          3948 => x"b8",
          3949 => x"d0",
          3950 => x"b8",
          3951 => x"ff",
          3952 => x"53",
          3953 => x"51",
          3954 => x"3f",
          3955 => x"d0",
          3956 => x"d0",
          3957 => x"57",
          3958 => x"2e",
          3959 => x"84",
          3960 => x"52",
          3961 => x"a7",
          3962 => x"d4",
          3963 => x"a0",
          3964 => x"fc",
          3965 => x"c8",
          3966 => x"51",
          3967 => x"3f",
          3968 => x"33",
          3969 => x"79",
          3970 => x"34",
          3971 => x"06",
          3972 => x"80",
          3973 => x"0b",
          3974 => x"34",
          3975 => x"d0",
          3976 => x"84",
          3977 => x"b4",
          3978 => x"75",
          3979 => x"fa",
          3980 => x"e4",
          3981 => x"a4",
          3982 => x"e4",
          3983 => x"06",
          3984 => x"75",
          3985 => x"ff",
          3986 => x"81",
          3987 => x"ff",
          3988 => x"a4",
          3989 => x"a8",
          3990 => x"5e",
          3991 => x"2e",
          3992 => x"84",
          3993 => x"52",
          3994 => x"a6",
          3995 => x"d4",
          3996 => x"a0",
          3997 => x"f8",
          3998 => x"c8",
          3999 => x"51",
          4000 => x"3f",
          4001 => x"33",
          4002 => x"76",
          4003 => x"34",
          4004 => x"06",
          4005 => x"75",
          4006 => x"8e",
          4007 => x"e4",
          4008 => x"a4",
          4009 => x"e4",
          4010 => x"06",
          4011 => x"75",
          4012 => x"ff",
          4013 => x"ff",
          4014 => x"ff",
          4015 => x"a4",
          4016 => x"a8",
          4017 => x"5e",
          4018 => x"2e",
          4019 => x"84",
          4020 => x"52",
          4021 => x"a5",
          4022 => x"d4",
          4023 => x"a0",
          4024 => x"8c",
          4025 => x"c8",
          4026 => x"51",
          4027 => x"3f",
          4028 => x"33",
          4029 => x"60",
          4030 => x"34",
          4031 => x"06",
          4032 => x"74",
          4033 => x"fa",
          4034 => x"d4",
          4035 => x"2b",
          4036 => x"83",
          4037 => x"81",
          4038 => x"52",
          4039 => x"dc",
          4040 => x"b8",
          4041 => x"0c",
          4042 => x"33",
          4043 => x"83",
          4044 => x"70",
          4045 => x"41",
          4046 => x"f4",
          4047 => x"53",
          4048 => x"51",
          4049 => x"3f",
          4050 => x"33",
          4051 => x"81",
          4052 => x"56",
          4053 => x"82",
          4054 => x"83",
          4055 => x"f4",
          4056 => x"3d",
          4057 => x"54",
          4058 => x"52",
          4059 => x"d8",
          4060 => x"f2",
          4061 => x"8a",
          4062 => x"88",
          4063 => x"d0",
          4064 => x"df",
          4065 => x"0b",
          4066 => x"34",
          4067 => x"d0",
          4068 => x"84",
          4069 => x"b4",
          4070 => x"93",
          4071 => x"84",
          4072 => x"51",
          4073 => x"3f",
          4074 => x"08",
          4075 => x"84",
          4076 => x"96",
          4077 => x"83",
          4078 => x"53",
          4079 => x"7a",
          4080 => x"f2",
          4081 => x"e4",
          4082 => x"b8",
          4083 => x"2e",
          4084 => x"e9",
          4085 => x"b8",
          4086 => x"ff",
          4087 => x"84",
          4088 => x"56",
          4089 => x"b8",
          4090 => x"80",
          4091 => x"b8",
          4092 => x"05",
          4093 => x"56",
          4094 => x"75",
          4095 => x"83",
          4096 => x"70",
          4097 => x"f1",
          4098 => x"08",
          4099 => x"59",
          4100 => x"38",
          4101 => x"87",
          4102 => x"f1",
          4103 => x"1a",
          4104 => x"55",
          4105 => x"3f",
          4106 => x"08",
          4107 => x"f2",
          4108 => x"10",
          4109 => x"fc",
          4110 => x"57",
          4111 => x"a0",
          4112 => x"70",
          4113 => x"5e",
          4114 => x"27",
          4115 => x"5d",
          4116 => x"09",
          4117 => x"df",
          4118 => x"ed",
          4119 => x"39",
          4120 => x"52",
          4121 => x"a6",
          4122 => x"f2",
          4123 => x"05",
          4124 => x"06",
          4125 => x"7a",
          4126 => x"38",
          4127 => x"f2",
          4128 => x"bd",
          4129 => x"80",
          4130 => x"83",
          4131 => x"70",
          4132 => x"fc",
          4133 => x"fc",
          4134 => x"70",
          4135 => x"57",
          4136 => x"3f",
          4137 => x"08",
          4138 => x"f2",
          4139 => x"10",
          4140 => x"fc",
          4141 => x"57",
          4142 => x"80",
          4143 => x"38",
          4144 => x"76",
          4145 => x"34",
          4146 => x"75",
          4147 => x"34",
          4148 => x"83",
          4149 => x"ff",
          4150 => x"77",
          4151 => x"f8",
          4152 => x"3d",
          4153 => x"c3",
          4154 => x"84",
          4155 => x"05",
          4156 => x"72",
          4157 => x"8d",
          4158 => x"2e",
          4159 => x"81",
          4160 => x"9e",
          4161 => x"2e",
          4162 => x"86",
          4163 => x"59",
          4164 => x"80",
          4165 => x"80",
          4166 => x"58",
          4167 => x"90",
          4168 => x"f8",
          4169 => x"83",
          4170 => x"75",
          4171 => x"23",
          4172 => x"33",
          4173 => x"71",
          4174 => x"71",
          4175 => x"71",
          4176 => x"56",
          4177 => x"78",
          4178 => x"38",
          4179 => x"84",
          4180 => x"74",
          4181 => x"05",
          4182 => x"74",
          4183 => x"75",
          4184 => x"38",
          4185 => x"33",
          4186 => x"17",
          4187 => x"55",
          4188 => x"0b",
          4189 => x"34",
          4190 => x"81",
          4191 => x"ff",
          4192 => x"ee",
          4193 => x"0d",
          4194 => x"a0",
          4195 => x"f8",
          4196 => x"10",
          4197 => x"f8",
          4198 => x"90",
          4199 => x"05",
          4200 => x"40",
          4201 => x"b0",
          4202 => x"b6",
          4203 => x"81",
          4204 => x"b6",
          4205 => x"81",
          4206 => x"f8",
          4207 => x"83",
          4208 => x"70",
          4209 => x"59",
          4210 => x"57",
          4211 => x"73",
          4212 => x"72",
          4213 => x"29",
          4214 => x"ff",
          4215 => x"ff",
          4216 => x"ff",
          4217 => x"ff",
          4218 => x"81",
          4219 => x"75",
          4220 => x"42",
          4221 => x"5c",
          4222 => x"8f",
          4223 => x"94",
          4224 => x"31",
          4225 => x"29",
          4226 => x"76",
          4227 => x"7b",
          4228 => x"9c",
          4229 => x"55",
          4230 => x"26",
          4231 => x"80",
          4232 => x"05",
          4233 => x"f8",
          4234 => x"70",
          4235 => x"34",
          4236 => x"a7",
          4237 => x"86",
          4238 => x"70",
          4239 => x"33",
          4240 => x"06",
          4241 => x"33",
          4242 => x"06",
          4243 => x"22",
          4244 => x"5d",
          4245 => x"5e",
          4246 => x"74",
          4247 => x"df",
          4248 => x"ff",
          4249 => x"ff",
          4250 => x"29",
          4251 => x"54",
          4252 => x"fd",
          4253 => x"0b",
          4254 => x"34",
          4255 => x"f8",
          4256 => x"f8",
          4257 => x"98",
          4258 => x"2b",
          4259 => x"2b",
          4260 => x"7a",
          4261 => x"56",
          4262 => x"26",
          4263 => x"fd",
          4264 => x"fc",
          4265 => x"f8",
          4266 => x"81",
          4267 => x"10",
          4268 => x"f8",
          4269 => x"90",
          4270 => x"a7",
          4271 => x"5e",
          4272 => x"56",
          4273 => x"b0",
          4274 => x"84",
          4275 => x"70",
          4276 => x"84",
          4277 => x"70",
          4278 => x"83",
          4279 => x"70",
          4280 => x"06",
          4281 => x"60",
          4282 => x"41",
          4283 => x"40",
          4284 => x"73",
          4285 => x"72",
          4286 => x"70",
          4287 => x"57",
          4288 => x"ff",
          4289 => x"ff",
          4290 => x"29",
          4291 => x"ff",
          4292 => x"ff",
          4293 => x"29",
          4294 => x"5c",
          4295 => x"78",
          4296 => x"77",
          4297 => x"79",
          4298 => x"79",
          4299 => x"58",
          4300 => x"38",
          4301 => x"5c",
          4302 => x"38",
          4303 => x"74",
          4304 => x"29",
          4305 => x"39",
          4306 => x"86",
          4307 => x"53",
          4308 => x"34",
          4309 => x"85",
          4310 => x"73",
          4311 => x"80",
          4312 => x"f4",
          4313 => x"b0",
          4314 => x"ee",
          4315 => x"80",
          4316 => x"76",
          4317 => x"80",
          4318 => x"74",
          4319 => x"34",
          4320 => x"34",
          4321 => x"51",
          4322 => x"86",
          4323 => x"70",
          4324 => x"81",
          4325 => x"a0",
          4326 => x"77",
          4327 => x"54",
          4328 => x"34",
          4329 => x"80",
          4330 => x"c0",
          4331 => x"72",
          4332 => x"a0",
          4333 => x"70",
          4334 => x"07",
          4335 => x"86",
          4336 => x"34",
          4337 => x"f7",
          4338 => x"53",
          4339 => x"80",
          4340 => x"b6",
          4341 => x"0b",
          4342 => x"0c",
          4343 => x"04",
          4344 => x"33",
          4345 => x"0c",
          4346 => x"0d",
          4347 => x"33",
          4348 => x"b3",
          4349 => x"b6",
          4350 => x"59",
          4351 => x"75",
          4352 => x"da",
          4353 => x"d8",
          4354 => x"95",
          4355 => x"94",
          4356 => x"29",
          4357 => x"a0",
          4358 => x"f8",
          4359 => x"51",
          4360 => x"7c",
          4361 => x"83",
          4362 => x"83",
          4363 => x"53",
          4364 => x"72",
          4365 => x"c4",
          4366 => x"92",
          4367 => x"55",
          4368 => x"92",
          4369 => x"94",
          4370 => x"70",
          4371 => x"7a",
          4372 => x"55",
          4373 => x"7a",
          4374 => x"38",
          4375 => x"72",
          4376 => x"34",
          4377 => x"22",
          4378 => x"ff",
          4379 => x"d6",
          4380 => x"57",
          4381 => x"82",
          4382 => x"b6",
          4383 => x"71",
          4384 => x"80",
          4385 => x"9f",
          4386 => x"84",
          4387 => x"14",
          4388 => x"e0",
          4389 => x"e0",
          4390 => x"70",
          4391 => x"33",
          4392 => x"05",
          4393 => x"14",
          4394 => x"d5",
          4395 => x"38",
          4396 => x"26",
          4397 => x"f8",
          4398 => x"97",
          4399 => x"55",
          4400 => x"e0",
          4401 => x"73",
          4402 => x"55",
          4403 => x"54",
          4404 => x"27",
          4405 => x"b6",
          4406 => x"05",
          4407 => x"f8",
          4408 => x"57",
          4409 => x"06",
          4410 => x"ff",
          4411 => x"73",
          4412 => x"fd",
          4413 => x"31",
          4414 => x"b6",
          4415 => x"71",
          4416 => x"57",
          4417 => x"a7",
          4418 => x"86",
          4419 => x"79",
          4420 => x"75",
          4421 => x"71",
          4422 => x"5c",
          4423 => x"75",
          4424 => x"38",
          4425 => x"16",
          4426 => x"14",
          4427 => x"b6",
          4428 => x"78",
          4429 => x"5a",
          4430 => x"81",
          4431 => x"77",
          4432 => x"59",
          4433 => x"84",
          4434 => x"84",
          4435 => x"71",
          4436 => x"56",
          4437 => x"72",
          4438 => x"38",
          4439 => x"84",
          4440 => x"8b",
          4441 => x"74",
          4442 => x"34",
          4443 => x"22",
          4444 => x"ff",
          4445 => x"d6",
          4446 => x"57",
          4447 => x"fd",
          4448 => x"80",
          4449 => x"38",
          4450 => x"06",
          4451 => x"f8",
          4452 => x"53",
          4453 => x"09",
          4454 => x"c8",
          4455 => x"31",
          4456 => x"b6",
          4457 => x"71",
          4458 => x"29",
          4459 => x"59",
          4460 => x"27",
          4461 => x"83",
          4462 => x"84",
          4463 => x"74",
          4464 => x"56",
          4465 => x"e0",
          4466 => x"75",
          4467 => x"05",
          4468 => x"13",
          4469 => x"2e",
          4470 => x"a0",
          4471 => x"16",
          4472 => x"70",
          4473 => x"34",
          4474 => x"72",
          4475 => x"f4",
          4476 => x"84",
          4477 => x"55",
          4478 => x"39",
          4479 => x"15",
          4480 => x"b6",
          4481 => x"74",
          4482 => x"d7",
          4483 => x"a9",
          4484 => x"0d",
          4485 => x"05",
          4486 => x"53",
          4487 => x"26",
          4488 => x"10",
          4489 => x"dc",
          4490 => x"08",
          4491 => x"d8",
          4492 => x"71",
          4493 => x"71",
          4494 => x"34",
          4495 => x"b8",
          4496 => x"3d",
          4497 => x"0b",
          4498 => x"34",
          4499 => x"33",
          4500 => x"06",
          4501 => x"80",
          4502 => x"ff",
          4503 => x"83",
          4504 => x"80",
          4505 => x"e4",
          4506 => x"0d",
          4507 => x"94",
          4508 => x"31",
          4509 => x"9f",
          4510 => x"54",
          4511 => x"70",
          4512 => x"34",
          4513 => x"f8",
          4514 => x"05",
          4515 => x"33",
          4516 => x"56",
          4517 => x"25",
          4518 => x"53",
          4519 => x"94",
          4520 => x"84",
          4521 => x"86",
          4522 => x"83",
          4523 => x"70",
          4524 => x"09",
          4525 => x"72",
          4526 => x"53",
          4527 => x"f8",
          4528 => x"0b",
          4529 => x"0c",
          4530 => x"04",
          4531 => x"33",
          4532 => x"b6",
          4533 => x"11",
          4534 => x"70",
          4535 => x"38",
          4536 => x"83",
          4537 => x"80",
          4538 => x"e4",
          4539 => x"0d",
          4540 => x"83",
          4541 => x"83",
          4542 => x"84",
          4543 => x"ff",
          4544 => x"71",
          4545 => x"b4",
          4546 => x"51",
          4547 => x"94",
          4548 => x"39",
          4549 => x"02",
          4550 => x"51",
          4551 => x"b3",
          4552 => x"10",
          4553 => x"05",
          4554 => x"04",
          4555 => x"33",
          4556 => x"06",
          4557 => x"80",
          4558 => x"72",
          4559 => x"51",
          4560 => x"71",
          4561 => x"09",
          4562 => x"38",
          4563 => x"83",
          4564 => x"80",
          4565 => x"e4",
          4566 => x"0d",
          4567 => x"90",
          4568 => x"06",
          4569 => x"70",
          4570 => x"34",
          4571 => x"b8",
          4572 => x"3d",
          4573 => x"f8",
          4574 => x"f0",
          4575 => x"83",
          4576 => x"e8",
          4577 => x"90",
          4578 => x"06",
          4579 => x"70",
          4580 => x"34",
          4581 => x"f1",
          4582 => x"90",
          4583 => x"84",
          4584 => x"83",
          4585 => x"83",
          4586 => x"81",
          4587 => x"07",
          4588 => x"f8",
          4589 => x"b4",
          4590 => x"90",
          4591 => x"51",
          4592 => x"90",
          4593 => x"39",
          4594 => x"33",
          4595 => x"85",
          4596 => x"83",
          4597 => x"ff",
          4598 => x"f8",
          4599 => x"fb",
          4600 => x"51",
          4601 => x"90",
          4602 => x"39",
          4603 => x"33",
          4604 => x"81",
          4605 => x"83",
          4606 => x"fe",
          4607 => x"f8",
          4608 => x"f8",
          4609 => x"83",
          4610 => x"fe",
          4611 => x"f8",
          4612 => x"df",
          4613 => x"07",
          4614 => x"f8",
          4615 => x"cc",
          4616 => x"90",
          4617 => x"06",
          4618 => x"70",
          4619 => x"34",
          4620 => x"83",
          4621 => x"81",
          4622 => x"e0",
          4623 => x"83",
          4624 => x"fe",
          4625 => x"f8",
          4626 => x"cf",
          4627 => x"07",
          4628 => x"f8",
          4629 => x"94",
          4630 => x"90",
          4631 => x"06",
          4632 => x"70",
          4633 => x"34",
          4634 => x"83",
          4635 => x"81",
          4636 => x"70",
          4637 => x"34",
          4638 => x"83",
          4639 => x"81",
          4640 => x"07",
          4641 => x"f8",
          4642 => x"e0",
          4643 => x"0d",
          4644 => x"33",
          4645 => x"80",
          4646 => x"83",
          4647 => x"83",
          4648 => x"83",
          4649 => x"84",
          4650 => x"43",
          4651 => x"5b",
          4652 => x"2e",
          4653 => x"78",
          4654 => x"38",
          4655 => x"81",
          4656 => x"84",
          4657 => x"80",
          4658 => x"dc",
          4659 => x"f8",
          4660 => x"83",
          4661 => x"7c",
          4662 => x"34",
          4663 => x"04",
          4664 => x"09",
          4665 => x"38",
          4666 => x"b6",
          4667 => x"0b",
          4668 => x"34",
          4669 => x"f8",
          4670 => x"0b",
          4671 => x"34",
          4672 => x"f8",
          4673 => x"58",
          4674 => x"33",
          4675 => x"d7",
          4676 => x"b6",
          4677 => x"7b",
          4678 => x"7a",
          4679 => x"d8",
          4680 => x"e6",
          4681 => x"b6",
          4682 => x"0b",
          4683 => x"34",
          4684 => x"94",
          4685 => x"f8",
          4686 => x"83",
          4687 => x"8f",
          4688 => x"80",
          4689 => x"da",
          4690 => x"84",
          4691 => x"80",
          4692 => x"94",
          4693 => x"83",
          4694 => x"80",
          4695 => x"92",
          4696 => x"e7",
          4697 => x"b7",
          4698 => x"84",
          4699 => x"56",
          4700 => x"54",
          4701 => x"52",
          4702 => x"51",
          4703 => x"3f",
          4704 => x"b7",
          4705 => x"5a",
          4706 => x"a5",
          4707 => x"84",
          4708 => x"70",
          4709 => x"83",
          4710 => x"ff",
          4711 => x"81",
          4712 => x"ff",
          4713 => x"e5",
          4714 => x"59",
          4715 => x"dd",
          4716 => x"94",
          4717 => x"d2",
          4718 => x"b6",
          4719 => x"0b",
          4720 => x"34",
          4721 => x"94",
          4722 => x"f8",
          4723 => x"83",
          4724 => x"8f",
          4725 => x"80",
          4726 => x"da",
          4727 => x"84",
          4728 => x"81",
          4729 => x"94",
          4730 => x"83",
          4731 => x"81",
          4732 => x"92",
          4733 => x"c8",
          4734 => x"ae",
          4735 => x"e4",
          4736 => x"e3",
          4737 => x"80",
          4738 => x"59",
          4739 => x"51",
          4740 => x"3f",
          4741 => x"e4",
          4742 => x"a6",
          4743 => x"c8",
          4744 => x"83",
          4745 => x"fe",
          4746 => x"81",
          4747 => x"ff",
          4748 => x"d8",
          4749 => x"0d",
          4750 => x"05",
          4751 => x"84",
          4752 => x"83",
          4753 => x"83",
          4754 => x"72",
          4755 => x"86",
          4756 => x"11",
          4757 => x"22",
          4758 => x"5c",
          4759 => x"05",
          4760 => x"ff",
          4761 => x"ea",
          4762 => x"51",
          4763 => x"72",
          4764 => x"e9",
          4765 => x"2e",
          4766 => x"75",
          4767 => x"b9",
          4768 => x"2e",
          4769 => x"75",
          4770 => x"d5",
          4771 => x"d8",
          4772 => x"94",
          4773 => x"95",
          4774 => x"29",
          4775 => x"54",
          4776 => x"16",
          4777 => x"a0",
          4778 => x"84",
          4779 => x"83",
          4780 => x"83",
          4781 => x"72",
          4782 => x"5a",
          4783 => x"75",
          4784 => x"18",
          4785 => x"94",
          4786 => x"29",
          4787 => x"83",
          4788 => x"86",
          4789 => x"18",
          4790 => x"d8",
          4791 => x"ff",
          4792 => x"92",
          4793 => x"95",
          4794 => x"29",
          4795 => x"57",
          4796 => x"f8",
          4797 => x"97",
          4798 => x"81",
          4799 => x"ff",
          4800 => x"73",
          4801 => x"99",
          4802 => x"d9",
          4803 => x"81",
          4804 => x"17",
          4805 => x"f8",
          4806 => x"b6",
          4807 => x"72",
          4808 => x"38",
          4809 => x"33",
          4810 => x"2e",
          4811 => x"80",
          4812 => x"e4",
          4813 => x"0d",
          4814 => x"2e",
          4815 => x"8d",
          4816 => x"38",
          4817 => x"09",
          4818 => x"c1",
          4819 => x"81",
          4820 => x"3f",
          4821 => x"f8",
          4822 => x"be",
          4823 => x"96",
          4824 => x"84",
          4825 => x"33",
          4826 => x"89",
          4827 => x"06",
          4828 => x"80",
          4829 => x"a0",
          4830 => x"3f",
          4831 => x"81",
          4832 => x"54",
          4833 => x"ff",
          4834 => x"52",
          4835 => x"a5",
          4836 => x"70",
          4837 => x"54",
          4838 => x"27",
          4839 => x"fa",
          4840 => x"f8",
          4841 => x"f2",
          4842 => x"83",
          4843 => x"3f",
          4844 => x"b8",
          4845 => x"3d",
          4846 => x"80",
          4847 => x"81",
          4848 => x"38",
          4849 => x"33",
          4850 => x"06",
          4851 => x"53",
          4852 => x"73",
          4853 => x"f8",
          4854 => x"52",
          4855 => x"d5",
          4856 => x"95",
          4857 => x"ff",
          4858 => x"05",
          4859 => x"a5",
          4860 => x"72",
          4861 => x"34",
          4862 => x"80",
          4863 => x"95",
          4864 => x"81",
          4865 => x"3f",
          4866 => x"80",
          4867 => x"ef",
          4868 => x"86",
          4869 => x"0d",
          4870 => x"05",
          4871 => x"e0",
          4872 => x"75",
          4873 => x"b8",
          4874 => x"2e",
          4875 => x"78",
          4876 => x"b5",
          4877 => x"24",
          4878 => x"78",
          4879 => x"b9",
          4880 => x"2e",
          4881 => x"84",
          4882 => x"83",
          4883 => x"83",
          4884 => x"72",
          4885 => x"58",
          4886 => x"b6",
          4887 => x"86",
          4888 => x"17",
          4889 => x"d8",
          4890 => x"95",
          4891 => x"92",
          4892 => x"29",
          4893 => x"42",
          4894 => x"f8",
          4895 => x"83",
          4896 => x"60",
          4897 => x"05",
          4898 => x"f8",
          4899 => x"86",
          4900 => x"05",
          4901 => x"d8",
          4902 => x"ff",
          4903 => x"92",
          4904 => x"95",
          4905 => x"29",
          4906 => x"5d",
          4907 => x"f8",
          4908 => x"97",
          4909 => x"81",
          4910 => x"ff",
          4911 => x"76",
          4912 => x"b8",
          4913 => x"d9",
          4914 => x"86",
          4915 => x"19",
          4916 => x"f8",
          4917 => x"0b",
          4918 => x"0c",
          4919 => x"04",
          4920 => x"84",
          4921 => x"79",
          4922 => x"38",
          4923 => x"9b",
          4924 => x"80",
          4925 => x"cc",
          4926 => x"84",
          4927 => x"84",
          4928 => x"83",
          4929 => x"83",
          4930 => x"72",
          4931 => x"5e",
          4932 => x"b6",
          4933 => x"86",
          4934 => x"1d",
          4935 => x"d8",
          4936 => x"95",
          4937 => x"92",
          4938 => x"29",
          4939 => x"59",
          4940 => x"f8",
          4941 => x"83",
          4942 => x"76",
          4943 => x"5b",
          4944 => x"90",
          4945 => x"b0",
          4946 => x"84",
          4947 => x"70",
          4948 => x"83",
          4949 => x"83",
          4950 => x"72",
          4951 => x"44",
          4952 => x"59",
          4953 => x"33",
          4954 => x"b6",
          4955 => x"1f",
          4956 => x"ff",
          4957 => x"77",
          4958 => x"38",
          4959 => x"95",
          4960 => x"84",
          4961 => x"9c",
          4962 => x"78",
          4963 => x"b7",
          4964 => x"24",
          4965 => x"78",
          4966 => x"81",
          4967 => x"38",
          4968 => x"f8",
          4969 => x"0b",
          4970 => x"0c",
          4971 => x"04",
          4972 => x"82",
          4973 => x"19",
          4974 => x"26",
          4975 => x"84",
          4976 => x"81",
          4977 => x"77",
          4978 => x"34",
          4979 => x"e8",
          4980 => x"81",
          4981 => x"80",
          4982 => x"e8",
          4983 => x"0b",
          4984 => x"0c",
          4985 => x"04",
          4986 => x"fd",
          4987 => x"0b",
          4988 => x"0c",
          4989 => x"33",
          4990 => x"33",
          4991 => x"33",
          4992 => x"05",
          4993 => x"84",
          4994 => x"33",
          4995 => x"80",
          4996 => x"b6",
          4997 => x"f8",
          4998 => x"f8",
          4999 => x"71",
          5000 => x"5f",
          5001 => x"83",
          5002 => x"34",
          5003 => x"33",
          5004 => x"19",
          5005 => x"f8",
          5006 => x"a7",
          5007 => x"34",
          5008 => x"33",
          5009 => x"06",
          5010 => x"22",
          5011 => x"33",
          5012 => x"11",
          5013 => x"58",
          5014 => x"90",
          5015 => x"97",
          5016 => x"81",
          5017 => x"89",
          5018 => x"81",
          5019 => x"3f",
          5020 => x"f8",
          5021 => x"ae",
          5022 => x"d8",
          5023 => x"95",
          5024 => x"ff",
          5025 => x"94",
          5026 => x"29",
          5027 => x"a0",
          5028 => x"f8",
          5029 => x"51",
          5030 => x"29",
          5031 => x"ff",
          5032 => x"f6",
          5033 => x"51",
          5034 => x"75",
          5035 => x"a4",
          5036 => x"ff",
          5037 => x"57",
          5038 => x"95",
          5039 => x"75",
          5040 => x"34",
          5041 => x"80",
          5042 => x"e4",
          5043 => x"84",
          5044 => x"80",
          5045 => x"e6",
          5046 => x"84",
          5047 => x"81",
          5048 => x"e0",
          5049 => x"84",
          5050 => x"9c",
          5051 => x"83",
          5052 => x"84",
          5053 => x"83",
          5054 => x"84",
          5055 => x"83",
          5056 => x"84",
          5057 => x"80",
          5058 => x"e0",
          5059 => x"84",
          5060 => x"9c",
          5061 => x"78",
          5062 => x"09",
          5063 => x"a7",
          5064 => x"94",
          5065 => x"d8",
          5066 => x"ff",
          5067 => x"95",
          5068 => x"ff",
          5069 => x"29",
          5070 => x"a0",
          5071 => x"f8",
          5072 => x"40",
          5073 => x"05",
          5074 => x"ff",
          5075 => x"ea",
          5076 => x"43",
          5077 => x"5c",
          5078 => x"85",
          5079 => x"81",
          5080 => x"1a",
          5081 => x"83",
          5082 => x"76",
          5083 => x"34",
          5084 => x"06",
          5085 => x"06",
          5086 => x"06",
          5087 => x"05",
          5088 => x"84",
          5089 => x"86",
          5090 => x"1e",
          5091 => x"d8",
          5092 => x"95",
          5093 => x"92",
          5094 => x"29",
          5095 => x"42",
          5096 => x"83",
          5097 => x"34",
          5098 => x"33",
          5099 => x"62",
          5100 => x"83",
          5101 => x"86",
          5102 => x"1a",
          5103 => x"d8",
          5104 => x"ff",
          5105 => x"92",
          5106 => x"95",
          5107 => x"29",
          5108 => x"5a",
          5109 => x"f8",
          5110 => x"84",
          5111 => x"34",
          5112 => x"81",
          5113 => x"58",
          5114 => x"95",
          5115 => x"b6",
          5116 => x"79",
          5117 => x"ff",
          5118 => x"83",
          5119 => x"83",
          5120 => x"70",
          5121 => x"58",
          5122 => x"fd",
          5123 => x"bb",
          5124 => x"38",
          5125 => x"83",
          5126 => x"bf",
          5127 => x"38",
          5128 => x"33",
          5129 => x"f9",
          5130 => x"19",
          5131 => x"26",
          5132 => x"75",
          5133 => x"c5",
          5134 => x"77",
          5135 => x"0b",
          5136 => x"34",
          5137 => x"51",
          5138 => x"80",
          5139 => x"e4",
          5140 => x"0d",
          5141 => x"94",
          5142 => x"d8",
          5143 => x"ff",
          5144 => x"95",
          5145 => x"ff",
          5146 => x"29",
          5147 => x"a0",
          5148 => x"f8",
          5149 => x"41",
          5150 => x"05",
          5151 => x"ff",
          5152 => x"ea",
          5153 => x"45",
          5154 => x"5b",
          5155 => x"82",
          5156 => x"5c",
          5157 => x"06",
          5158 => x"06",
          5159 => x"06",
          5160 => x"05",
          5161 => x"84",
          5162 => x"86",
          5163 => x"1b",
          5164 => x"d8",
          5165 => x"95",
          5166 => x"92",
          5167 => x"29",
          5168 => x"5e",
          5169 => x"83",
          5170 => x"34",
          5171 => x"33",
          5172 => x"1e",
          5173 => x"f8",
          5174 => x"a7",
          5175 => x"34",
          5176 => x"33",
          5177 => x"06",
          5178 => x"22",
          5179 => x"33",
          5180 => x"11",
          5181 => x"40",
          5182 => x"90",
          5183 => x"b6",
          5184 => x"81",
          5185 => x"ff",
          5186 => x"7e",
          5187 => x"ac",
          5188 => x"d9",
          5189 => x"92",
          5190 => x"19",
          5191 => x"f8",
          5192 => x"1c",
          5193 => x"06",
          5194 => x"83",
          5195 => x"38",
          5196 => x"33",
          5197 => x"33",
          5198 => x"33",
          5199 => x"06",
          5200 => x"06",
          5201 => x"06",
          5202 => x"05",
          5203 => x"5b",
          5204 => x"b7",
          5205 => x"a7",
          5206 => x"34",
          5207 => x"33",
          5208 => x"33",
          5209 => x"22",
          5210 => x"12",
          5211 => x"56",
          5212 => x"f8",
          5213 => x"83",
          5214 => x"76",
          5215 => x"5a",
          5216 => x"90",
          5217 => x"b0",
          5218 => x"84",
          5219 => x"70",
          5220 => x"83",
          5221 => x"83",
          5222 => x"72",
          5223 => x"5b",
          5224 => x"59",
          5225 => x"33",
          5226 => x"18",
          5227 => x"05",
          5228 => x"06",
          5229 => x"7f",
          5230 => x"38",
          5231 => x"95",
          5232 => x"39",
          5233 => x"b7",
          5234 => x"0b",
          5235 => x"0c",
          5236 => x"04",
          5237 => x"17",
          5238 => x"b6",
          5239 => x"7a",
          5240 => x"95",
          5241 => x"ff",
          5242 => x"05",
          5243 => x"39",
          5244 => x"b7",
          5245 => x"0b",
          5246 => x"0c",
          5247 => x"04",
          5248 => x"17",
          5249 => x"b6",
          5250 => x"7c",
          5251 => x"94",
          5252 => x"d8",
          5253 => x"95",
          5254 => x"5b",
          5255 => x"f4",
          5256 => x"e8",
          5257 => x"dc",
          5258 => x"05",
          5259 => x"d8",
          5260 => x"e4",
          5261 => x"fb",
          5262 => x"b7",
          5263 => x"11",
          5264 => x"84",
          5265 => x"79",
          5266 => x"06",
          5267 => x"ca",
          5268 => x"84",
          5269 => x"23",
          5270 => x"83",
          5271 => x"33",
          5272 => x"e0",
          5273 => x"34",
          5274 => x"33",
          5275 => x"33",
          5276 => x"33",
          5277 => x"f9",
          5278 => x"b6",
          5279 => x"f8",
          5280 => x"f8",
          5281 => x"72",
          5282 => x"5d",
          5283 => x"e0",
          5284 => x"86",
          5285 => x"05",
          5286 => x"d8",
          5287 => x"95",
          5288 => x"92",
          5289 => x"29",
          5290 => x"5b",
          5291 => x"f8",
          5292 => x"83",
          5293 => x"76",
          5294 => x"41",
          5295 => x"90",
          5296 => x"a7",
          5297 => x"34",
          5298 => x"33",
          5299 => x"06",
          5300 => x"22",
          5301 => x"33",
          5302 => x"11",
          5303 => x"42",
          5304 => x"90",
          5305 => x"b6",
          5306 => x"1c",
          5307 => x"06",
          5308 => x"7b",
          5309 => x"38",
          5310 => x"33",
          5311 => x"e2",
          5312 => x"56",
          5313 => x"95",
          5314 => x"84",
          5315 => x"84",
          5316 => x"40",
          5317 => x"f3",
          5318 => x"b6",
          5319 => x"75",
          5320 => x"78",
          5321 => x"ea",
          5322 => x"0b",
          5323 => x"0c",
          5324 => x"04",
          5325 => x"33",
          5326 => x"34",
          5327 => x"33",
          5328 => x"34",
          5329 => x"33",
          5330 => x"f8",
          5331 => x"b9",
          5332 => x"94",
          5333 => x"cc",
          5334 => x"95",
          5335 => x"cd",
          5336 => x"93",
          5337 => x"ce",
          5338 => x"39",
          5339 => x"33",
          5340 => x"2e",
          5341 => x"84",
          5342 => x"5d",
          5343 => x"09",
          5344 => x"85",
          5345 => x"95",
          5346 => x"55",
          5347 => x"33",
          5348 => x"9b",
          5349 => x"a0",
          5350 => x"70",
          5351 => x"ee",
          5352 => x"51",
          5353 => x"3f",
          5354 => x"08",
          5355 => x"83",
          5356 => x"57",
          5357 => x"60",
          5358 => x"cd",
          5359 => x"83",
          5360 => x"fe",
          5361 => x"fe",
          5362 => x"0b",
          5363 => x"33",
          5364 => x"81",
          5365 => x"77",
          5366 => x"ad",
          5367 => x"84",
          5368 => x"81",
          5369 => x"41",
          5370 => x"8a",
          5371 => x"10",
          5372 => x"94",
          5373 => x"08",
          5374 => x"e5",
          5375 => x"80",
          5376 => x"38",
          5377 => x"33",
          5378 => x"33",
          5379 => x"70",
          5380 => x"2c",
          5381 => x"42",
          5382 => x"75",
          5383 => x"34",
          5384 => x"84",
          5385 => x"56",
          5386 => x"8e",
          5387 => x"b8",
          5388 => x"05",
          5389 => x"06",
          5390 => x"33",
          5391 => x"75",
          5392 => x"c5",
          5393 => x"f8",
          5394 => x"bd",
          5395 => x"83",
          5396 => x"83",
          5397 => x"70",
          5398 => x"5d",
          5399 => x"2e",
          5400 => x"ff",
          5401 => x"83",
          5402 => x"fd",
          5403 => x"0b",
          5404 => x"34",
          5405 => x"33",
          5406 => x"33",
          5407 => x"57",
          5408 => x"fd",
          5409 => x"17",
          5410 => x"f8",
          5411 => x"f9",
          5412 => x"e5",
          5413 => x"80",
          5414 => x"38",
          5415 => x"33",
          5416 => x"33",
          5417 => x"70",
          5418 => x"2c",
          5419 => x"41",
          5420 => x"75",
          5421 => x"34",
          5422 => x"84",
          5423 => x"5b",
          5424 => x"fc",
          5425 => x"b8",
          5426 => x"60",
          5427 => x"81",
          5428 => x"38",
          5429 => x"33",
          5430 => x"33",
          5431 => x"33",
          5432 => x"12",
          5433 => x"80",
          5434 => x"92",
          5435 => x"5a",
          5436 => x"29",
          5437 => x"ff",
          5438 => x"f6",
          5439 => x"ff",
          5440 => x"42",
          5441 => x"7e",
          5442 => x"2e",
          5443 => x"80",
          5444 => x"e9",
          5445 => x"39",
          5446 => x"33",
          5447 => x"2e",
          5448 => x"84",
          5449 => x"58",
          5450 => x"09",
          5451 => x"d9",
          5452 => x"83",
          5453 => x"fb",
          5454 => x"b7",
          5455 => x"75",
          5456 => x"be",
          5457 => x"b9",
          5458 => x"95",
          5459 => x"05",
          5460 => x"33",
          5461 => x"5e",
          5462 => x"25",
          5463 => x"57",
          5464 => x"95",
          5465 => x"39",
          5466 => x"33",
          5467 => x"2e",
          5468 => x"84",
          5469 => x"83",
          5470 => x"42",
          5471 => x"b6",
          5472 => x"11",
          5473 => x"75",
          5474 => x"38",
          5475 => x"83",
          5476 => x"fa",
          5477 => x"e3",
          5478 => x"e8",
          5479 => x"0b",
          5480 => x"33",
          5481 => x"76",
          5482 => x"38",
          5483 => x"b8",
          5484 => x"22",
          5485 => x"e3",
          5486 => x"e8",
          5487 => x"17",
          5488 => x"06",
          5489 => x"33",
          5490 => x"da",
          5491 => x"84",
          5492 => x"5f",
          5493 => x"2e",
          5494 => x"b8",
          5495 => x"75",
          5496 => x"38",
          5497 => x"52",
          5498 => x"06",
          5499 => x"3f",
          5500 => x"84",
          5501 => x"57",
          5502 => x"8e",
          5503 => x"b8",
          5504 => x"05",
          5505 => x"06",
          5506 => x"33",
          5507 => x"81",
          5508 => x"b6",
          5509 => x"81",
          5510 => x"11",
          5511 => x"5b",
          5512 => x"77",
          5513 => x"38",
          5514 => x"83",
          5515 => x"76",
          5516 => x"ff",
          5517 => x"77",
          5518 => x"38",
          5519 => x"83",
          5520 => x"84",
          5521 => x"ff",
          5522 => x"7a",
          5523 => x"b4",
          5524 => x"75",
          5525 => x"34",
          5526 => x"84",
          5527 => x"5f",
          5528 => x"8a",
          5529 => x"b8",
          5530 => x"b6",
          5531 => x"5b",
          5532 => x"f9",
          5533 => x"f8",
          5534 => x"b6",
          5535 => x"81",
          5536 => x"f8",
          5537 => x"74",
          5538 => x"a7",
          5539 => x"83",
          5540 => x"5f",
          5541 => x"29",
          5542 => x"ff",
          5543 => x"f6",
          5544 => x"52",
          5545 => x"5d",
          5546 => x"84",
          5547 => x"83",
          5548 => x"70",
          5549 => x"57",
          5550 => x"8e",
          5551 => x"b6",
          5552 => x"76",
          5553 => x"d6",
          5554 => x"56",
          5555 => x"92",
          5556 => x"ff",
          5557 => x"31",
          5558 => x"60",
          5559 => x"38",
          5560 => x"33",
          5561 => x"27",
          5562 => x"ff",
          5563 => x"83",
          5564 => x"7e",
          5565 => x"83",
          5566 => x"57",
          5567 => x"76",
          5568 => x"38",
          5569 => x"81",
          5570 => x"ff",
          5571 => x"29",
          5572 => x"79",
          5573 => x"a0",
          5574 => x"a7",
          5575 => x"81",
          5576 => x"81",
          5577 => x"71",
          5578 => x"58",
          5579 => x"7f",
          5580 => x"38",
          5581 => x"1a",
          5582 => x"17",
          5583 => x"b6",
          5584 => x"7b",
          5585 => x"5d",
          5586 => x"81",
          5587 => x"7c",
          5588 => x"5e",
          5589 => x"84",
          5590 => x"84",
          5591 => x"71",
          5592 => x"43",
          5593 => x"77",
          5594 => x"9d",
          5595 => x"17",
          5596 => x"b6",
          5597 => x"7b",
          5598 => x"5d",
          5599 => x"81",
          5600 => x"7c",
          5601 => x"5e",
          5602 => x"84",
          5603 => x"84",
          5604 => x"71",
          5605 => x"43",
          5606 => x"7f",
          5607 => x"99",
          5608 => x"39",
          5609 => x"33",
          5610 => x"2e",
          5611 => x"80",
          5612 => x"b9",
          5613 => x"b1",
          5614 => x"39",
          5615 => x"b6",
          5616 => x"11",
          5617 => x"33",
          5618 => x"58",
          5619 => x"94",
          5620 => x"b8",
          5621 => x"78",
          5622 => x"06",
          5623 => x"83",
          5624 => x"58",
          5625 => x"06",
          5626 => x"33",
          5627 => x"5c",
          5628 => x"81",
          5629 => x"b6",
          5630 => x"7a",
          5631 => x"89",
          5632 => x"ff",
          5633 => x"76",
          5634 => x"38",
          5635 => x"61",
          5636 => x"57",
          5637 => x"38",
          5638 => x"1b",
          5639 => x"62",
          5640 => x"a0",
          5641 => x"1f",
          5642 => x"a7",
          5643 => x"79",
          5644 => x"51",
          5645 => x"ac",
          5646 => x"06",
          5647 => x"a4",
          5648 => x"90",
          5649 => x"2b",
          5650 => x"07",
          5651 => x"07",
          5652 => x"7f",
          5653 => x"57",
          5654 => x"9e",
          5655 => x"70",
          5656 => x"0c",
          5657 => x"84",
          5658 => x"79",
          5659 => x"38",
          5660 => x"33",
          5661 => x"33",
          5662 => x"81",
          5663 => x"81",
          5664 => x"f8",
          5665 => x"73",
          5666 => x"59",
          5667 => x"77",
          5668 => x"38",
          5669 => x"1b",
          5670 => x"62",
          5671 => x"75",
          5672 => x"57",
          5673 => x"f4",
          5674 => x"f8",
          5675 => x"97",
          5676 => x"5a",
          5677 => x"e0",
          5678 => x"78",
          5679 => x"5a",
          5680 => x"57",
          5681 => x"f4",
          5682 => x"0b",
          5683 => x"34",
          5684 => x"81",
          5685 => x"81",
          5686 => x"77",
          5687 => x"f4",
          5688 => x"1f",
          5689 => x"06",
          5690 => x"8a",
          5691 => x"90",
          5692 => x"f0",
          5693 => x"2b",
          5694 => x"71",
          5695 => x"58",
          5696 => x"80",
          5697 => x"81",
          5698 => x"80",
          5699 => x"f8",
          5700 => x"18",
          5701 => x"06",
          5702 => x"b6",
          5703 => x"96",
          5704 => x"84",
          5705 => x"33",
          5706 => x"f8",
          5707 => x"b6",
          5708 => x"f8",
          5709 => x"b6",
          5710 => x"5c",
          5711 => x"ee",
          5712 => x"90",
          5713 => x"56",
          5714 => x"90",
          5715 => x"70",
          5716 => x"59",
          5717 => x"39",
          5718 => x"33",
          5719 => x"85",
          5720 => x"83",
          5721 => x"e5",
          5722 => x"90",
          5723 => x"06",
          5724 => x"75",
          5725 => x"34",
          5726 => x"f8",
          5727 => x"f9",
          5728 => x"56",
          5729 => x"90",
          5730 => x"83",
          5731 => x"81",
          5732 => x"07",
          5733 => x"f8",
          5734 => x"b1",
          5735 => x"0b",
          5736 => x"34",
          5737 => x"81",
          5738 => x"56",
          5739 => x"83",
          5740 => x"81",
          5741 => x"75",
          5742 => x"34",
          5743 => x"83",
          5744 => x"81",
          5745 => x"07",
          5746 => x"f8",
          5747 => x"fd",
          5748 => x"90",
          5749 => x"06",
          5750 => x"56",
          5751 => x"90",
          5752 => x"39",
          5753 => x"33",
          5754 => x"80",
          5755 => x"75",
          5756 => x"34",
          5757 => x"83",
          5758 => x"81",
          5759 => x"07",
          5760 => x"f8",
          5761 => x"c5",
          5762 => x"90",
          5763 => x"06",
          5764 => x"75",
          5765 => x"34",
          5766 => x"83",
          5767 => x"81",
          5768 => x"07",
          5769 => x"f8",
          5770 => x"a1",
          5771 => x"90",
          5772 => x"06",
          5773 => x"75",
          5774 => x"34",
          5775 => x"83",
          5776 => x"81",
          5777 => x"75",
          5778 => x"34",
          5779 => x"83",
          5780 => x"80",
          5781 => x"75",
          5782 => x"34",
          5783 => x"83",
          5784 => x"80",
          5785 => x"75",
          5786 => x"34",
          5787 => x"83",
          5788 => x"81",
          5789 => x"d0",
          5790 => x"83",
          5791 => x"fd",
          5792 => x"f8",
          5793 => x"bf",
          5794 => x"56",
          5795 => x"90",
          5796 => x"39",
          5797 => x"f8",
          5798 => x"52",
          5799 => x"c9",
          5800 => x"39",
          5801 => x"33",
          5802 => x"34",
          5803 => x"33",
          5804 => x"34",
          5805 => x"33",
          5806 => x"f8",
          5807 => x"0b",
          5808 => x"0c",
          5809 => x"81",
          5810 => x"e7",
          5811 => x"84",
          5812 => x"9c",
          5813 => x"77",
          5814 => x"34",
          5815 => x"33",
          5816 => x"06",
          5817 => x"56",
          5818 => x"84",
          5819 => x"9c",
          5820 => x"53",
          5821 => x"fe",
          5822 => x"84",
          5823 => x"a1",
          5824 => x"e4",
          5825 => x"e0",
          5826 => x"84",
          5827 => x"80",
          5828 => x"e4",
          5829 => x"0d",
          5830 => x"f8",
          5831 => x"e9",
          5832 => x"e5",
          5833 => x"5c",
          5834 => x"b7",
          5835 => x"10",
          5836 => x"5d",
          5837 => x"05",
          5838 => x"b8",
          5839 => x"0b",
          5840 => x"34",
          5841 => x"0b",
          5842 => x"34",
          5843 => x"51",
          5844 => x"83",
          5845 => x"70",
          5846 => x"58",
          5847 => x"e6",
          5848 => x"0b",
          5849 => x"34",
          5850 => x"51",
          5851 => x"ef",
          5852 => x"51",
          5853 => x"3f",
          5854 => x"83",
          5855 => x"ff",
          5856 => x"70",
          5857 => x"06",
          5858 => x"f2",
          5859 => x"52",
          5860 => x"39",
          5861 => x"33",
          5862 => x"27",
          5863 => x"75",
          5864 => x"34",
          5865 => x"83",
          5866 => x"ff",
          5867 => x"70",
          5868 => x"06",
          5869 => x"f0",
          5870 => x"f8",
          5871 => x"05",
          5872 => x"33",
          5873 => x"59",
          5874 => x"25",
          5875 => x"75",
          5876 => x"39",
          5877 => x"33",
          5878 => x"06",
          5879 => x"77",
          5880 => x"38",
          5881 => x"33",
          5882 => x"33",
          5883 => x"06",
          5884 => x"33",
          5885 => x"11",
          5886 => x"80",
          5887 => x"92",
          5888 => x"71",
          5889 => x"70",
          5890 => x"06",
          5891 => x"33",
          5892 => x"42",
          5893 => x"81",
          5894 => x"38",
          5895 => x"ff",
          5896 => x"5c",
          5897 => x"24",
          5898 => x"84",
          5899 => x"56",
          5900 => x"83",
          5901 => x"16",
          5902 => x"f8",
          5903 => x"81",
          5904 => x"11",
          5905 => x"76",
          5906 => x"38",
          5907 => x"33",
          5908 => x"27",
          5909 => x"ff",
          5910 => x"83",
          5911 => x"7b",
          5912 => x"83",
          5913 => x"57",
          5914 => x"76",
          5915 => x"38",
          5916 => x"81",
          5917 => x"ff",
          5918 => x"29",
          5919 => x"79",
          5920 => x"a0",
          5921 => x"a7",
          5922 => x"81",
          5923 => x"81",
          5924 => x"71",
          5925 => x"42",
          5926 => x"7e",
          5927 => x"38",
          5928 => x"1a",
          5929 => x"17",
          5930 => x"b6",
          5931 => x"7b",
          5932 => x"5d",
          5933 => x"81",
          5934 => x"7d",
          5935 => x"5f",
          5936 => x"84",
          5937 => x"84",
          5938 => x"71",
          5939 => x"59",
          5940 => x"77",
          5941 => x"b1",
          5942 => x"17",
          5943 => x"b6",
          5944 => x"7b",
          5945 => x"5d",
          5946 => x"81",
          5947 => x"7d",
          5948 => x"5f",
          5949 => x"84",
          5950 => x"84",
          5951 => x"71",
          5952 => x"59",
          5953 => x"75",
          5954 => x"99",
          5955 => x"39",
          5956 => x"17",
          5957 => x"b6",
          5958 => x"7b",
          5959 => x"94",
          5960 => x"d8",
          5961 => x"92",
          5962 => x"d7",
          5963 => x"5f",
          5964 => x"39",
          5965 => x"38",
          5966 => x"33",
          5967 => x"06",
          5968 => x"42",
          5969 => x"27",
          5970 => x"5a",
          5971 => x"92",
          5972 => x"ff",
          5973 => x"58",
          5974 => x"27",
          5975 => x"57",
          5976 => x"94",
          5977 => x"d8",
          5978 => x"ff",
          5979 => x"52",
          5980 => x"78",
          5981 => x"38",
          5982 => x"83",
          5983 => x"eb",
          5984 => x"f8",
          5985 => x"05",
          5986 => x"33",
          5987 => x"40",
          5988 => x"25",
          5989 => x"75",
          5990 => x"39",
          5991 => x"09",
          5992 => x"c0",
          5993 => x"95",
          5994 => x"ff",
          5995 => x"94",
          5996 => x"5d",
          5997 => x"ff",
          5998 => x"06",
          5999 => x"f6",
          6000 => x"1d",
          6001 => x"f8",
          6002 => x"93",
          6003 => x"56",
          6004 => x"92",
          6005 => x"39",
          6006 => x"56",
          6007 => x"94",
          6008 => x"39",
          6009 => x"56",
          6010 => x"f5",
          6011 => x"76",
          6012 => x"58",
          6013 => x"90",
          6014 => x"81",
          6015 => x"75",
          6016 => x"ec",
          6017 => x"70",
          6018 => x"34",
          6019 => x"33",
          6020 => x"05",
          6021 => x"76",
          6022 => x"f4",
          6023 => x"7b",
          6024 => x"83",
          6025 => x"f1",
          6026 => x"0b",
          6027 => x"34",
          6028 => x"7e",
          6029 => x"23",
          6030 => x"80",
          6031 => x"92",
          6032 => x"39",
          6033 => x"f8",
          6034 => x"a7",
          6035 => x"96",
          6036 => x"84",
          6037 => x"33",
          6038 => x"0b",
          6039 => x"34",
          6040 => x"fd",
          6041 => x"97",
          6042 => x"b6",
          6043 => x"54",
          6044 => x"90",
          6045 => x"db",
          6046 => x"0b",
          6047 => x"0c",
          6048 => x"04",
          6049 => x"51",
          6050 => x"80",
          6051 => x"e4",
          6052 => x"0d",
          6053 => x"0d",
          6054 => x"33",
          6055 => x"83",
          6056 => x"70",
          6057 => x"83",
          6058 => x"33",
          6059 => x"59",
          6060 => x"80",
          6061 => x"14",
          6062 => x"f6",
          6063 => x"59",
          6064 => x"e4",
          6065 => x"0d",
          6066 => x"c4",
          6067 => x"53",
          6068 => x"91",
          6069 => x"32",
          6070 => x"07",
          6071 => x"9f",
          6072 => x"5e",
          6073 => x"f6",
          6074 => x"59",
          6075 => x"81",
          6076 => x"06",
          6077 => x"54",
          6078 => x"70",
          6079 => x"25",
          6080 => x"5c",
          6081 => x"2e",
          6082 => x"84",
          6083 => x"83",
          6084 => x"83",
          6085 => x"72",
          6086 => x"86",
          6087 => x"05",
          6088 => x"22",
          6089 => x"71",
          6090 => x"70",
          6091 => x"06",
          6092 => x"33",
          6093 => x"58",
          6094 => x"83",
          6095 => x"f0",
          6096 => x"ee",
          6097 => x"80",
          6098 => x"98",
          6099 => x"c0",
          6100 => x"56",
          6101 => x"f6",
          6102 => x"80",
          6103 => x"76",
          6104 => x"15",
          6105 => x"70",
          6106 => x"55",
          6107 => x"74",
          6108 => x"80",
          6109 => x"84",
          6110 => x"81",
          6111 => x"f6",
          6112 => x"58",
          6113 => x"76",
          6114 => x"38",
          6115 => x"2e",
          6116 => x"74",
          6117 => x"15",
          6118 => x"ff",
          6119 => x"81",
          6120 => x"cd",
          6121 => x"f6",
          6122 => x"83",
          6123 => x"33",
          6124 => x"15",
          6125 => x"70",
          6126 => x"55",
          6127 => x"27",
          6128 => x"83",
          6129 => x"70",
          6130 => x"80",
          6131 => x"54",
          6132 => x"bc",
          6133 => x"ff",
          6134 => x"2a",
          6135 => x"81",
          6136 => x"58",
          6137 => x"85",
          6138 => x"0b",
          6139 => x"34",
          6140 => x"06",
          6141 => x"2e",
          6142 => x"81",
          6143 => x"be",
          6144 => x"83",
          6145 => x"83",
          6146 => x"83",
          6147 => x"70",
          6148 => x"33",
          6149 => x"33",
          6150 => x"5e",
          6151 => x"83",
          6152 => x"33",
          6153 => x"ff",
          6154 => x"83",
          6155 => x"33",
          6156 => x"2e",
          6157 => x"83",
          6158 => x"33",
          6159 => x"ff",
          6160 => x"83",
          6161 => x"33",
          6162 => x"ec",
          6163 => x"ff",
          6164 => x"81",
          6165 => x"38",
          6166 => x"16",
          6167 => x"81",
          6168 => x"38",
          6169 => x"06",
          6170 => x"ff",
          6171 => x"38",
          6172 => x"16",
          6173 => x"74",
          6174 => x"38",
          6175 => x"08",
          6176 => x"87",
          6177 => x"08",
          6178 => x"73",
          6179 => x"38",
          6180 => x"c0",
          6181 => x"83",
          6182 => x"58",
          6183 => x"81",
          6184 => x"54",
          6185 => x"fe",
          6186 => x"83",
          6187 => x"77",
          6188 => x"34",
          6189 => x"53",
          6190 => x"82",
          6191 => x"10",
          6192 => x"dc",
          6193 => x"08",
          6194 => x"ec",
          6195 => x"80",
          6196 => x"83",
          6197 => x"c0",
          6198 => x"5e",
          6199 => x"27",
          6200 => x"80",
          6201 => x"ea",
          6202 => x"72",
          6203 => x"38",
          6204 => x"83",
          6205 => x"87",
          6206 => x"08",
          6207 => x"0c",
          6208 => x"06",
          6209 => x"2e",
          6210 => x"f8",
          6211 => x"54",
          6212 => x"14",
          6213 => x"81",
          6214 => x"a5",
          6215 => x"c4",
          6216 => x"80",
          6217 => x"38",
          6218 => x"83",
          6219 => x"c3",
          6220 => x"f0",
          6221 => x"39",
          6222 => x"e0",
          6223 => x"56",
          6224 => x"7c",
          6225 => x"38",
          6226 => x"09",
          6227 => x"b4",
          6228 => x"2e",
          6229 => x"79",
          6230 => x"d7",
          6231 => x"ff",
          6232 => x"77",
          6233 => x"2b",
          6234 => x"80",
          6235 => x"73",
          6236 => x"38",
          6237 => x"81",
          6238 => x"10",
          6239 => x"87",
          6240 => x"98",
          6241 => x"57",
          6242 => x"73",
          6243 => x"78",
          6244 => x"79",
          6245 => x"11",
          6246 => x"05",
          6247 => x"05",
          6248 => x"56",
          6249 => x"c0",
          6250 => x"83",
          6251 => x"57",
          6252 => x"80",
          6253 => x"2e",
          6254 => x"79",
          6255 => x"59",
          6256 => x"82",
          6257 => x"39",
          6258 => x"fa",
          6259 => x"0b",
          6260 => x"33",
          6261 => x"81",
          6262 => x"38",
          6263 => x"70",
          6264 => x"25",
          6265 => x"59",
          6266 => x"38",
          6267 => x"09",
          6268 => x"cc",
          6269 => x"2e",
          6270 => x"80",
          6271 => x"10",
          6272 => x"f0",
          6273 => x"5d",
          6274 => x"2e",
          6275 => x"81",
          6276 => x"ff",
          6277 => x"93",
          6278 => x"38",
          6279 => x"33",
          6280 => x"2e",
          6281 => x"84",
          6282 => x"55",
          6283 => x"38",
          6284 => x"06",
          6285 => x"cc",
          6286 => x"84",
          6287 => x"8f",
          6288 => x"be",
          6289 => x"f0",
          6290 => x"39",
          6291 => x"2e",
          6292 => x"f6",
          6293 => x"81",
          6294 => x"83",
          6295 => x"34",
          6296 => x"80",
          6297 => x"ac",
          6298 => x"0b",
          6299 => x"15",
          6300 => x"83",
          6301 => x"34",
          6302 => x"74",
          6303 => x"53",
          6304 => x"2e",
          6305 => x"83",
          6306 => x"33",
          6307 => x"27",
          6308 => x"77",
          6309 => x"54",
          6310 => x"09",
          6311 => x"fc",
          6312 => x"b8",
          6313 => x"05",
          6314 => x"9c",
          6315 => x"74",
          6316 => x"e8",
          6317 => x"98",
          6318 => x"f6",
          6319 => x"81",
          6320 => x"fb",
          6321 => x"0b",
          6322 => x"15",
          6323 => x"39",
          6324 => x"bd",
          6325 => x"81",
          6326 => x"fa",
          6327 => x"83",
          6328 => x"80",
          6329 => x"bd",
          6330 => x"c4",
          6331 => x"be",
          6332 => x"f6",
          6333 => x"f6",
          6334 => x"5d",
          6335 => x"5e",
          6336 => x"39",
          6337 => x"09",
          6338 => x"cb",
          6339 => x"7a",
          6340 => x"ce",
          6341 => x"2e",
          6342 => x"fc",
          6343 => x"93",
          6344 => x"34",
          6345 => x"f8",
          6346 => x"0b",
          6347 => x"33",
          6348 => x"83",
          6349 => x"73",
          6350 => x"34",
          6351 => x"ac",
          6352 => x"84",
          6353 => x"58",
          6354 => x"38",
          6355 => x"84",
          6356 => x"ff",
          6357 => x"39",
          6358 => x"f6",
          6359 => x"2e",
          6360 => x"84",
          6361 => x"c4",
          6362 => x"39",
          6363 => x"33",
          6364 => x"06",
          6365 => x"5a",
          6366 => x"27",
          6367 => x"55",
          6368 => x"92",
          6369 => x"ff",
          6370 => x"55",
          6371 => x"27",
          6372 => x"54",
          6373 => x"94",
          6374 => x"d8",
          6375 => x"ff",
          6376 => x"05",
          6377 => x"27",
          6378 => x"53",
          6379 => x"95",
          6380 => x"f6",
          6381 => x"52",
          6382 => x"ba",
          6383 => x"59",
          6384 => x"72",
          6385 => x"39",
          6386 => x"52",
          6387 => x"51",
          6388 => x"3f",
          6389 => x"f6",
          6390 => x"f6",
          6391 => x"fc",
          6392 => x"3d",
          6393 => x"f5",
          6394 => x"3d",
          6395 => x"3d",
          6396 => x"83",
          6397 => x"53",
          6398 => x"05",
          6399 => x"34",
          6400 => x"08",
          6401 => x"71",
          6402 => x"83",
          6403 => x"55",
          6404 => x"81",
          6405 => x"0b",
          6406 => x"e8",
          6407 => x"98",
          6408 => x"f2",
          6409 => x"80",
          6410 => x"53",
          6411 => x"9c",
          6412 => x"c0",
          6413 => x"51",
          6414 => x"f6",
          6415 => x"33",
          6416 => x"9c",
          6417 => x"74",
          6418 => x"38",
          6419 => x"2e",
          6420 => x"c0",
          6421 => x"51",
          6422 => x"73",
          6423 => x"38",
          6424 => x"ff",
          6425 => x"38",
          6426 => x"9c",
          6427 => x"90",
          6428 => x"c0",
          6429 => x"52",
          6430 => x"9c",
          6431 => x"72",
          6432 => x"81",
          6433 => x"c0",
          6434 => x"52",
          6435 => x"27",
          6436 => x"81",
          6437 => x"38",
          6438 => x"a4",
          6439 => x"75",
          6440 => x"ff",
          6441 => x"ff",
          6442 => x"ff",
          6443 => x"75",
          6444 => x"38",
          6445 => x"06",
          6446 => x"d5",
          6447 => x"2e",
          6448 => x"84",
          6449 => x"88",
          6450 => x"81",
          6451 => x"e4",
          6452 => x"0d",
          6453 => x"0d",
          6454 => x"05",
          6455 => x"56",
          6456 => x"83",
          6457 => x"73",
          6458 => x"fc",
          6459 => x"70",
          6460 => x"07",
          6461 => x"57",
          6462 => x"34",
          6463 => x"51",
          6464 => x"34",
          6465 => x"56",
          6466 => x"34",
          6467 => x"34",
          6468 => x"08",
          6469 => x"13",
          6470 => x"f0",
          6471 => x"e1",
          6472 => x"0b",
          6473 => x"08",
          6474 => x"0b",
          6475 => x"80",
          6476 => x"80",
          6477 => x"c0",
          6478 => x"83",
          6479 => x"55",
          6480 => x"05",
          6481 => x"98",
          6482 => x"87",
          6483 => x"08",
          6484 => x"2e",
          6485 => x"14",
          6486 => x"98",
          6487 => x"52",
          6488 => x"87",
          6489 => x"fe",
          6490 => x"87",
          6491 => x"08",
          6492 => x"70",
          6493 => x"c8",
          6494 => x"71",
          6495 => x"c0",
          6496 => x"98",
          6497 => x"ce",
          6498 => x"87",
          6499 => x"08",
          6500 => x"98",
          6501 => x"74",
          6502 => x"38",
          6503 => x"87",
          6504 => x"08",
          6505 => x"73",
          6506 => x"71",
          6507 => x"db",
          6508 => x"98",
          6509 => x"72",
          6510 => x"38",
          6511 => x"55",
          6512 => x"81",
          6513 => x"53",
          6514 => x"80",
          6515 => x"81",
          6516 => x"71",
          6517 => x"74",
          6518 => x"ff",
          6519 => x"aa",
          6520 => x"14",
          6521 => x"11",
          6522 => x"70",
          6523 => x"38",
          6524 => x"05",
          6525 => x"70",
          6526 => x"34",
          6527 => x"f0",
          6528 => x"b8",
          6529 => x"3d",
          6530 => x"0b",
          6531 => x"0c",
          6532 => x"04",
          6533 => x"39",
          6534 => x"79",
          6535 => x"a3",
          6536 => x"56",
          6537 => x"f2",
          6538 => x"88",
          6539 => x"80",
          6540 => x"79",
          6541 => x"51",
          6542 => x"75",
          6543 => x"72",
          6544 => x"70",
          6545 => x"75",
          6546 => x"71",
          6547 => x"72",
          6548 => x"7a",
          6549 => x"08",
          6550 => x"84",
          6551 => x"54",
          6552 => x"73",
          6553 => x"70",
          6554 => x"52",
          6555 => x"81",
          6556 => x"72",
          6557 => x"38",
          6558 => x"08",
          6559 => x"15",
          6560 => x"f0",
          6561 => x"e2",
          6562 => x"0b",
          6563 => x"08",
          6564 => x"0b",
          6565 => x"80",
          6566 => x"80",
          6567 => x"c0",
          6568 => x"83",
          6569 => x"55",
          6570 => x"05",
          6571 => x"98",
          6572 => x"87",
          6573 => x"08",
          6574 => x"2e",
          6575 => x"14",
          6576 => x"98",
          6577 => x"52",
          6578 => x"87",
          6579 => x"fe",
          6580 => x"87",
          6581 => x"08",
          6582 => x"70",
          6583 => x"c8",
          6584 => x"71",
          6585 => x"c0",
          6586 => x"98",
          6587 => x"ce",
          6588 => x"87",
          6589 => x"08",
          6590 => x"98",
          6591 => x"74",
          6592 => x"38",
          6593 => x"87",
          6594 => x"08",
          6595 => x"73",
          6596 => x"71",
          6597 => x"db",
          6598 => x"98",
          6599 => x"72",
          6600 => x"38",
          6601 => x"55",
          6602 => x"81",
          6603 => x"53",
          6604 => x"a1",
          6605 => x"ff",
          6606 => x"fe",
          6607 => x"51",
          6608 => x"06",
          6609 => x"2e",
          6610 => x"57",
          6611 => x"e4",
          6612 => x"0d",
          6613 => x"e8",
          6614 => x"0d",
          6615 => x"08",
          6616 => x"71",
          6617 => x"83",
          6618 => x"56",
          6619 => x"81",
          6620 => x"0b",
          6621 => x"e8",
          6622 => x"98",
          6623 => x"f2",
          6624 => x"80",
          6625 => x"54",
          6626 => x"9c",
          6627 => x"c0",
          6628 => x"53",
          6629 => x"f6",
          6630 => x"33",
          6631 => x"9c",
          6632 => x"70",
          6633 => x"38",
          6634 => x"2e",
          6635 => x"c0",
          6636 => x"51",
          6637 => x"74",
          6638 => x"38",
          6639 => x"ff",
          6640 => x"38",
          6641 => x"9c",
          6642 => x"90",
          6643 => x"c0",
          6644 => x"52",
          6645 => x"9c",
          6646 => x"72",
          6647 => x"81",
          6648 => x"c0",
          6649 => x"55",
          6650 => x"27",
          6651 => x"81",
          6652 => x"38",
          6653 => x"a4",
          6654 => x"71",
          6655 => x"ff",
          6656 => x"ff",
          6657 => x"ff",
          6658 => x"75",
          6659 => x"38",
          6660 => x"06",
          6661 => x"d5",
          6662 => x"80",
          6663 => x"e3",
          6664 => x"d0",
          6665 => x"3d",
          6666 => x"3d",
          6667 => x"d4",
          6668 => x"31",
          6669 => x"83",
          6670 => x"70",
          6671 => x"11",
          6672 => x"12",
          6673 => x"2b",
          6674 => x"07",
          6675 => x"33",
          6676 => x"71",
          6677 => x"90",
          6678 => x"54",
          6679 => x"5d",
          6680 => x"56",
          6681 => x"71",
          6682 => x"38",
          6683 => x"11",
          6684 => x"33",
          6685 => x"71",
          6686 => x"76",
          6687 => x"81",
          6688 => x"98",
          6689 => x"2b",
          6690 => x"5c",
          6691 => x"52",
          6692 => x"83",
          6693 => x"13",
          6694 => x"33",
          6695 => x"71",
          6696 => x"75",
          6697 => x"2a",
          6698 => x"57",
          6699 => x"34",
          6700 => x"06",
          6701 => x"13",
          6702 => x"d4",
          6703 => x"84",
          6704 => x"13",
          6705 => x"2b",
          6706 => x"2a",
          6707 => x"54",
          6708 => x"14",
          6709 => x"14",
          6710 => x"d4",
          6711 => x"80",
          6712 => x"34",
          6713 => x"13",
          6714 => x"d4",
          6715 => x"84",
          6716 => x"85",
          6717 => x"b8",
          6718 => x"70",
          6719 => x"33",
          6720 => x"07",
          6721 => x"07",
          6722 => x"58",
          6723 => x"74",
          6724 => x"81",
          6725 => x"3d",
          6726 => x"12",
          6727 => x"33",
          6728 => x"71",
          6729 => x"75",
          6730 => x"33",
          6731 => x"71",
          6732 => x"70",
          6733 => x"58",
          6734 => x"58",
          6735 => x"12",
          6736 => x"12",
          6737 => x"d4",
          6738 => x"84",
          6739 => x"12",
          6740 => x"2b",
          6741 => x"07",
          6742 => x"52",
          6743 => x"12",
          6744 => x"33",
          6745 => x"07",
          6746 => x"52",
          6747 => x"77",
          6748 => x"72",
          6749 => x"84",
          6750 => x"15",
          6751 => x"12",
          6752 => x"2b",
          6753 => x"ff",
          6754 => x"2a",
          6755 => x"52",
          6756 => x"77",
          6757 => x"84",
          6758 => x"70",
          6759 => x"81",
          6760 => x"8b",
          6761 => x"2b",
          6762 => x"70",
          6763 => x"33",
          6764 => x"07",
          6765 => x"8f",
          6766 => x"77",
          6767 => x"2a",
          6768 => x"54",
          6769 => x"54",
          6770 => x"14",
          6771 => x"14",
          6772 => x"d4",
          6773 => x"70",
          6774 => x"33",
          6775 => x"71",
          6776 => x"74",
          6777 => x"81",
          6778 => x"88",
          6779 => x"ff",
          6780 => x"88",
          6781 => x"53",
          6782 => x"54",
          6783 => x"34",
          6784 => x"34",
          6785 => x"08",
          6786 => x"11",
          6787 => x"33",
          6788 => x"71",
          6789 => x"74",
          6790 => x"81",
          6791 => x"98",
          6792 => x"2b",
          6793 => x"5d",
          6794 => x"53",
          6795 => x"25",
          6796 => x"71",
          6797 => x"33",
          6798 => x"07",
          6799 => x"07",
          6800 => x"59",
          6801 => x"75",
          6802 => x"16",
          6803 => x"d4",
          6804 => x"70",
          6805 => x"33",
          6806 => x"71",
          6807 => x"74",
          6808 => x"33",
          6809 => x"71",
          6810 => x"70",
          6811 => x"5c",
          6812 => x"56",
          6813 => x"82",
          6814 => x"83",
          6815 => x"3d",
          6816 => x"3d",
          6817 => x"b8",
          6818 => x"58",
          6819 => x"8f",
          6820 => x"2e",
          6821 => x"51",
          6822 => x"89",
          6823 => x"84",
          6824 => x"84",
          6825 => x"a0",
          6826 => x"b8",
          6827 => x"80",
          6828 => x"52",
          6829 => x"51",
          6830 => x"3f",
          6831 => x"08",
          6832 => x"34",
          6833 => x"16",
          6834 => x"d4",
          6835 => x"84",
          6836 => x"0b",
          6837 => x"84",
          6838 => x"56",
          6839 => x"34",
          6840 => x"17",
          6841 => x"d4",
          6842 => x"d0",
          6843 => x"fe",
          6844 => x"70",
          6845 => x"06",
          6846 => x"58",
          6847 => x"74",
          6848 => x"73",
          6849 => x"84",
          6850 => x"70",
          6851 => x"84",
          6852 => x"05",
          6853 => x"55",
          6854 => x"34",
          6855 => x"15",
          6856 => x"39",
          6857 => x"7b",
          6858 => x"81",
          6859 => x"27",
          6860 => x"12",
          6861 => x"05",
          6862 => x"ff",
          6863 => x"70",
          6864 => x"06",
          6865 => x"08",
          6866 => x"85",
          6867 => x"88",
          6868 => x"52",
          6869 => x"55",
          6870 => x"54",
          6871 => x"80",
          6872 => x"10",
          6873 => x"70",
          6874 => x"33",
          6875 => x"07",
          6876 => x"ff",
          6877 => x"70",
          6878 => x"06",
          6879 => x"56",
          6880 => x"54",
          6881 => x"27",
          6882 => x"80",
          6883 => x"75",
          6884 => x"84",
          6885 => x"13",
          6886 => x"2b",
          6887 => x"75",
          6888 => x"81",
          6889 => x"85",
          6890 => x"54",
          6891 => x"83",
          6892 => x"70",
          6893 => x"33",
          6894 => x"07",
          6895 => x"ff",
          6896 => x"5d",
          6897 => x"70",
          6898 => x"38",
          6899 => x"51",
          6900 => x"82",
          6901 => x"51",
          6902 => x"82",
          6903 => x"75",
          6904 => x"38",
          6905 => x"83",
          6906 => x"74",
          6907 => x"07",
          6908 => x"5b",
          6909 => x"5a",
          6910 => x"78",
          6911 => x"84",
          6912 => x"15",
          6913 => x"53",
          6914 => x"14",
          6915 => x"14",
          6916 => x"d4",
          6917 => x"70",
          6918 => x"33",
          6919 => x"07",
          6920 => x"8f",
          6921 => x"74",
          6922 => x"ff",
          6923 => x"88",
          6924 => x"53",
          6925 => x"52",
          6926 => x"34",
          6927 => x"06",
          6928 => x"12",
          6929 => x"d4",
          6930 => x"75",
          6931 => x"81",
          6932 => x"b8",
          6933 => x"19",
          6934 => x"87",
          6935 => x"8b",
          6936 => x"2b",
          6937 => x"58",
          6938 => x"57",
          6939 => x"34",
          6940 => x"34",
          6941 => x"08",
          6942 => x"78",
          6943 => x"33",
          6944 => x"71",
          6945 => x"70",
          6946 => x"54",
          6947 => x"86",
          6948 => x"87",
          6949 => x"b8",
          6950 => x"19",
          6951 => x"85",
          6952 => x"8b",
          6953 => x"2b",
          6954 => x"58",
          6955 => x"52",
          6956 => x"34",
          6957 => x"34",
          6958 => x"08",
          6959 => x"78",
          6960 => x"33",
          6961 => x"71",
          6962 => x"70",
          6963 => x"5c",
          6964 => x"84",
          6965 => x"85",
          6966 => x"b8",
          6967 => x"84",
          6968 => x"84",
          6969 => x"8b",
          6970 => x"86",
          6971 => x"15",
          6972 => x"2b",
          6973 => x"07",
          6974 => x"17",
          6975 => x"33",
          6976 => x"07",
          6977 => x"5a",
          6978 => x"54",
          6979 => x"12",
          6980 => x"12",
          6981 => x"d4",
          6982 => x"84",
          6983 => x"12",
          6984 => x"2b",
          6985 => x"07",
          6986 => x"14",
          6987 => x"33",
          6988 => x"07",
          6989 => x"58",
          6990 => x"56",
          6991 => x"70",
          6992 => x"76",
          6993 => x"84",
          6994 => x"18",
          6995 => x"12",
          6996 => x"2b",
          6997 => x"ff",
          6998 => x"2a",
          6999 => x"57",
          7000 => x"74",
          7001 => x"84",
          7002 => x"18",
          7003 => x"fe",
          7004 => x"3d",
          7005 => x"b8",
          7006 => x"58",
          7007 => x"a0",
          7008 => x"77",
          7009 => x"84",
          7010 => x"89",
          7011 => x"77",
          7012 => x"3f",
          7013 => x"08",
          7014 => x"0c",
          7015 => x"04",
          7016 => x"0b",
          7017 => x"0c",
          7018 => x"84",
          7019 => x"82",
          7020 => x"76",
          7021 => x"f4",
          7022 => x"c5",
          7023 => x"d4",
          7024 => x"75",
          7025 => x"81",
          7026 => x"b8",
          7027 => x"76",
          7028 => x"81",
          7029 => x"34",
          7030 => x"08",
          7031 => x"17",
          7032 => x"87",
          7033 => x"b8",
          7034 => x"b8",
          7035 => x"05",
          7036 => x"07",
          7037 => x"ff",
          7038 => x"2a",
          7039 => x"56",
          7040 => x"34",
          7041 => x"34",
          7042 => x"22",
          7043 => x"10",
          7044 => x"08",
          7045 => x"55",
          7046 => x"15",
          7047 => x"83",
          7048 => x"54",
          7049 => x"fe",
          7050 => x"e3",
          7051 => x"0d",
          7052 => x"5f",
          7053 => x"b8",
          7054 => x"45",
          7055 => x"2e",
          7056 => x"7e",
          7057 => x"af",
          7058 => x"2e",
          7059 => x"81",
          7060 => x"27",
          7061 => x"fb",
          7062 => x"82",
          7063 => x"ff",
          7064 => x"58",
          7065 => x"ff",
          7066 => x"31",
          7067 => x"83",
          7068 => x"70",
          7069 => x"11",
          7070 => x"12",
          7071 => x"2b",
          7072 => x"31",
          7073 => x"ff",
          7074 => x"10",
          7075 => x"73",
          7076 => x"11",
          7077 => x"12",
          7078 => x"2b",
          7079 => x"2b",
          7080 => x"53",
          7081 => x"44",
          7082 => x"44",
          7083 => x"52",
          7084 => x"80",
          7085 => x"fd",
          7086 => x"33",
          7087 => x"71",
          7088 => x"70",
          7089 => x"19",
          7090 => x"12",
          7091 => x"2b",
          7092 => x"07",
          7093 => x"56",
          7094 => x"74",
          7095 => x"38",
          7096 => x"82",
          7097 => x"1b",
          7098 => x"2e",
          7099 => x"60",
          7100 => x"f9",
          7101 => x"58",
          7102 => x"87",
          7103 => x"18",
          7104 => x"24",
          7105 => x"76",
          7106 => x"81",
          7107 => x"8b",
          7108 => x"2b",
          7109 => x"70",
          7110 => x"33",
          7111 => x"71",
          7112 => x"47",
          7113 => x"53",
          7114 => x"80",
          7115 => x"ba",
          7116 => x"82",
          7117 => x"12",
          7118 => x"2b",
          7119 => x"07",
          7120 => x"11",
          7121 => x"33",
          7122 => x"71",
          7123 => x"7e",
          7124 => x"33",
          7125 => x"71",
          7126 => x"70",
          7127 => x"57",
          7128 => x"41",
          7129 => x"59",
          7130 => x"1d",
          7131 => x"1d",
          7132 => x"d4",
          7133 => x"84",
          7134 => x"12",
          7135 => x"2b",
          7136 => x"07",
          7137 => x"14",
          7138 => x"33",
          7139 => x"07",
          7140 => x"5f",
          7141 => x"40",
          7142 => x"77",
          7143 => x"7b",
          7144 => x"84",
          7145 => x"16",
          7146 => x"12",
          7147 => x"2b",
          7148 => x"ff",
          7149 => x"2a",
          7150 => x"59",
          7151 => x"79",
          7152 => x"84",
          7153 => x"70",
          7154 => x"33",
          7155 => x"71",
          7156 => x"83",
          7157 => x"05",
          7158 => x"15",
          7159 => x"2b",
          7160 => x"2a",
          7161 => x"5d",
          7162 => x"55",
          7163 => x"75",
          7164 => x"84",
          7165 => x"70",
          7166 => x"81",
          7167 => x"8b",
          7168 => x"2b",
          7169 => x"82",
          7170 => x"15",
          7171 => x"2b",
          7172 => x"2a",
          7173 => x"5d",
          7174 => x"55",
          7175 => x"34",
          7176 => x"34",
          7177 => x"08",
          7178 => x"11",
          7179 => x"33",
          7180 => x"07",
          7181 => x"56",
          7182 => x"42",
          7183 => x"7e",
          7184 => x"51",
          7185 => x"3f",
          7186 => x"08",
          7187 => x"61",
          7188 => x"70",
          7189 => x"06",
          7190 => x"7a",
          7191 => x"b6",
          7192 => x"73",
          7193 => x"0c",
          7194 => x"04",
          7195 => x"0b",
          7196 => x"0c",
          7197 => x"84",
          7198 => x"82",
          7199 => x"60",
          7200 => x"f4",
          7201 => x"f9",
          7202 => x"d4",
          7203 => x"7e",
          7204 => x"81",
          7205 => x"b8",
          7206 => x"60",
          7207 => x"81",
          7208 => x"34",
          7209 => x"08",
          7210 => x"1d",
          7211 => x"87",
          7212 => x"b8",
          7213 => x"b8",
          7214 => x"05",
          7215 => x"07",
          7216 => x"ff",
          7217 => x"2a",
          7218 => x"57",
          7219 => x"34",
          7220 => x"34",
          7221 => x"22",
          7222 => x"10",
          7223 => x"08",
          7224 => x"55",
          7225 => x"15",
          7226 => x"83",
          7227 => x"b8",
          7228 => x"7e",
          7229 => x"76",
          7230 => x"8c",
          7231 => x"7f",
          7232 => x"df",
          7233 => x"f4",
          7234 => x"b8",
          7235 => x"b8",
          7236 => x"3d",
          7237 => x"1c",
          7238 => x"08",
          7239 => x"71",
          7240 => x"7f",
          7241 => x"81",
          7242 => x"88",
          7243 => x"ff",
          7244 => x"88",
          7245 => x"5b",
          7246 => x"7b",
          7247 => x"1c",
          7248 => x"b8",
          7249 => x"7c",
          7250 => x"58",
          7251 => x"34",
          7252 => x"34",
          7253 => x"08",
          7254 => x"33",
          7255 => x"71",
          7256 => x"70",
          7257 => x"ff",
          7258 => x"05",
          7259 => x"ff",
          7260 => x"2a",
          7261 => x"57",
          7262 => x"63",
          7263 => x"34",
          7264 => x"06",
          7265 => x"83",
          7266 => x"b8",
          7267 => x"5b",
          7268 => x"60",
          7269 => x"61",
          7270 => x"08",
          7271 => x"51",
          7272 => x"7e",
          7273 => x"39",
          7274 => x"70",
          7275 => x"06",
          7276 => x"ac",
          7277 => x"ff",
          7278 => x"31",
          7279 => x"ff",
          7280 => x"33",
          7281 => x"71",
          7282 => x"70",
          7283 => x"1b",
          7284 => x"12",
          7285 => x"2b",
          7286 => x"07",
          7287 => x"54",
          7288 => x"54",
          7289 => x"f9",
          7290 => x"bc",
          7291 => x"24",
          7292 => x"80",
          7293 => x"8f",
          7294 => x"ff",
          7295 => x"61",
          7296 => x"dd",
          7297 => x"39",
          7298 => x"0b",
          7299 => x"0c",
          7300 => x"84",
          7301 => x"82",
          7302 => x"7e",
          7303 => x"f4",
          7304 => x"dd",
          7305 => x"d4",
          7306 => x"7a",
          7307 => x"81",
          7308 => x"b8",
          7309 => x"7e",
          7310 => x"81",
          7311 => x"34",
          7312 => x"08",
          7313 => x"19",
          7314 => x"87",
          7315 => x"b8",
          7316 => x"b8",
          7317 => x"05",
          7318 => x"07",
          7319 => x"ff",
          7320 => x"2a",
          7321 => x"44",
          7322 => x"05",
          7323 => x"89",
          7324 => x"b8",
          7325 => x"10",
          7326 => x"b8",
          7327 => x"f8",
          7328 => x"7e",
          7329 => x"34",
          7330 => x"05",
          7331 => x"39",
          7332 => x"83",
          7333 => x"83",
          7334 => x"5b",
          7335 => x"fb",
          7336 => x"f2",
          7337 => x"2e",
          7338 => x"7e",
          7339 => x"3f",
          7340 => x"84",
          7341 => x"95",
          7342 => x"76",
          7343 => x"33",
          7344 => x"71",
          7345 => x"83",
          7346 => x"11",
          7347 => x"87",
          7348 => x"8b",
          7349 => x"2b",
          7350 => x"84",
          7351 => x"15",
          7352 => x"2b",
          7353 => x"2a",
          7354 => x"56",
          7355 => x"53",
          7356 => x"78",
          7357 => x"34",
          7358 => x"05",
          7359 => x"d4",
          7360 => x"84",
          7361 => x"12",
          7362 => x"2b",
          7363 => x"07",
          7364 => x"14",
          7365 => x"33",
          7366 => x"07",
          7367 => x"5b",
          7368 => x"5d",
          7369 => x"73",
          7370 => x"34",
          7371 => x"05",
          7372 => x"d4",
          7373 => x"33",
          7374 => x"71",
          7375 => x"81",
          7376 => x"70",
          7377 => x"5c",
          7378 => x"7d",
          7379 => x"1e",
          7380 => x"d4",
          7381 => x"82",
          7382 => x"12",
          7383 => x"2b",
          7384 => x"07",
          7385 => x"33",
          7386 => x"71",
          7387 => x"70",
          7388 => x"5c",
          7389 => x"57",
          7390 => x"7c",
          7391 => x"1d",
          7392 => x"d4",
          7393 => x"70",
          7394 => x"33",
          7395 => x"71",
          7396 => x"74",
          7397 => x"33",
          7398 => x"71",
          7399 => x"70",
          7400 => x"47",
          7401 => x"5c",
          7402 => x"82",
          7403 => x"83",
          7404 => x"b8",
          7405 => x"1f",
          7406 => x"83",
          7407 => x"88",
          7408 => x"57",
          7409 => x"83",
          7410 => x"58",
          7411 => x"84",
          7412 => x"bd",
          7413 => x"b8",
          7414 => x"84",
          7415 => x"ff",
          7416 => x"5f",
          7417 => x"84",
          7418 => x"84",
          7419 => x"a0",
          7420 => x"b8",
          7421 => x"80",
          7422 => x"52",
          7423 => x"51",
          7424 => x"3f",
          7425 => x"08",
          7426 => x"34",
          7427 => x"17",
          7428 => x"d4",
          7429 => x"84",
          7430 => x"0b",
          7431 => x"84",
          7432 => x"54",
          7433 => x"34",
          7434 => x"15",
          7435 => x"d4",
          7436 => x"d0",
          7437 => x"fe",
          7438 => x"70",
          7439 => x"06",
          7440 => x"45",
          7441 => x"61",
          7442 => x"60",
          7443 => x"84",
          7444 => x"70",
          7445 => x"84",
          7446 => x"05",
          7447 => x"5d",
          7448 => x"34",
          7449 => x"1c",
          7450 => x"e7",
          7451 => x"54",
          7452 => x"86",
          7453 => x"1a",
          7454 => x"2b",
          7455 => x"07",
          7456 => x"1c",
          7457 => x"33",
          7458 => x"07",
          7459 => x"5c",
          7460 => x"59",
          7461 => x"84",
          7462 => x"61",
          7463 => x"84",
          7464 => x"70",
          7465 => x"33",
          7466 => x"71",
          7467 => x"83",
          7468 => x"05",
          7469 => x"87",
          7470 => x"88",
          7471 => x"88",
          7472 => x"48",
          7473 => x"59",
          7474 => x"86",
          7475 => x"64",
          7476 => x"84",
          7477 => x"1d",
          7478 => x"12",
          7479 => x"2b",
          7480 => x"ff",
          7481 => x"2a",
          7482 => x"58",
          7483 => x"7f",
          7484 => x"84",
          7485 => x"70",
          7486 => x"81",
          7487 => x"8b",
          7488 => x"2b",
          7489 => x"70",
          7490 => x"33",
          7491 => x"07",
          7492 => x"8f",
          7493 => x"77",
          7494 => x"2a",
          7495 => x"5a",
          7496 => x"44",
          7497 => x"17",
          7498 => x"17",
          7499 => x"d4",
          7500 => x"70",
          7501 => x"33",
          7502 => x"71",
          7503 => x"74",
          7504 => x"81",
          7505 => x"88",
          7506 => x"ff",
          7507 => x"88",
          7508 => x"5e",
          7509 => x"41",
          7510 => x"34",
          7511 => x"05",
          7512 => x"ff",
          7513 => x"fa",
          7514 => x"15",
          7515 => x"33",
          7516 => x"71",
          7517 => x"79",
          7518 => x"33",
          7519 => x"71",
          7520 => x"70",
          7521 => x"5e",
          7522 => x"5d",
          7523 => x"34",
          7524 => x"34",
          7525 => x"08",
          7526 => x"11",
          7527 => x"33",
          7528 => x"71",
          7529 => x"74",
          7530 => x"33",
          7531 => x"71",
          7532 => x"70",
          7533 => x"56",
          7534 => x"42",
          7535 => x"60",
          7536 => x"75",
          7537 => x"34",
          7538 => x"08",
          7539 => x"81",
          7540 => x"88",
          7541 => x"ff",
          7542 => x"88",
          7543 => x"58",
          7544 => x"34",
          7545 => x"34",
          7546 => x"08",
          7547 => x"33",
          7548 => x"71",
          7549 => x"83",
          7550 => x"05",
          7551 => x"12",
          7552 => x"2b",
          7553 => x"2b",
          7554 => x"06",
          7555 => x"88",
          7556 => x"5f",
          7557 => x"42",
          7558 => x"82",
          7559 => x"83",
          7560 => x"b8",
          7561 => x"1f",
          7562 => x"12",
          7563 => x"2b",
          7564 => x"07",
          7565 => x"33",
          7566 => x"71",
          7567 => x"81",
          7568 => x"70",
          7569 => x"54",
          7570 => x"59",
          7571 => x"7c",
          7572 => x"1d",
          7573 => x"d4",
          7574 => x"82",
          7575 => x"12",
          7576 => x"2b",
          7577 => x"07",
          7578 => x"11",
          7579 => x"33",
          7580 => x"71",
          7581 => x"78",
          7582 => x"33",
          7583 => x"71",
          7584 => x"70",
          7585 => x"57",
          7586 => x"42",
          7587 => x"5a",
          7588 => x"84",
          7589 => x"85",
          7590 => x"b8",
          7591 => x"17",
          7592 => x"85",
          7593 => x"8b",
          7594 => x"2b",
          7595 => x"86",
          7596 => x"15",
          7597 => x"2b",
          7598 => x"2a",
          7599 => x"52",
          7600 => x"57",
          7601 => x"34",
          7602 => x"34",
          7603 => x"08",
          7604 => x"81",
          7605 => x"88",
          7606 => x"ff",
          7607 => x"88",
          7608 => x"5e",
          7609 => x"34",
          7610 => x"34",
          7611 => x"08",
          7612 => x"11",
          7613 => x"33",
          7614 => x"71",
          7615 => x"74",
          7616 => x"81",
          7617 => x"88",
          7618 => x"88",
          7619 => x"45",
          7620 => x"55",
          7621 => x"34",
          7622 => x"34",
          7623 => x"08",
          7624 => x"33",
          7625 => x"71",
          7626 => x"83",
          7627 => x"05",
          7628 => x"83",
          7629 => x"88",
          7630 => x"88",
          7631 => x"45",
          7632 => x"55",
          7633 => x"1a",
          7634 => x"1a",
          7635 => x"d4",
          7636 => x"82",
          7637 => x"12",
          7638 => x"2b",
          7639 => x"62",
          7640 => x"2b",
          7641 => x"5d",
          7642 => x"05",
          7643 => x"d4",
          7644 => x"d4",
          7645 => x"05",
          7646 => x"1c",
          7647 => x"ff",
          7648 => x"5f",
          7649 => x"86",
          7650 => x"1a",
          7651 => x"2b",
          7652 => x"07",
          7653 => x"1c",
          7654 => x"33",
          7655 => x"07",
          7656 => x"40",
          7657 => x"41",
          7658 => x"84",
          7659 => x"61",
          7660 => x"84",
          7661 => x"70",
          7662 => x"33",
          7663 => x"71",
          7664 => x"83",
          7665 => x"05",
          7666 => x"87",
          7667 => x"88",
          7668 => x"88",
          7669 => x"5f",
          7670 => x"41",
          7671 => x"86",
          7672 => x"64",
          7673 => x"84",
          7674 => x"1d",
          7675 => x"12",
          7676 => x"2b",
          7677 => x"ff",
          7678 => x"2a",
          7679 => x"55",
          7680 => x"7c",
          7681 => x"84",
          7682 => x"70",
          7683 => x"81",
          7684 => x"8b",
          7685 => x"2b",
          7686 => x"70",
          7687 => x"33",
          7688 => x"07",
          7689 => x"8f",
          7690 => x"77",
          7691 => x"2a",
          7692 => x"49",
          7693 => x"58",
          7694 => x"1e",
          7695 => x"1e",
          7696 => x"d4",
          7697 => x"70",
          7698 => x"33",
          7699 => x"71",
          7700 => x"74",
          7701 => x"81",
          7702 => x"88",
          7703 => x"ff",
          7704 => x"88",
          7705 => x"49",
          7706 => x"5e",
          7707 => x"34",
          7708 => x"34",
          7709 => x"ff",
          7710 => x"83",
          7711 => x"52",
          7712 => x"3f",
          7713 => x"08",
          7714 => x"e4",
          7715 => x"93",
          7716 => x"73",
          7717 => x"e4",
          7718 => x"b5",
          7719 => x"51",
          7720 => x"61",
          7721 => x"27",
          7722 => x"f0",
          7723 => x"3d",
          7724 => x"29",
          7725 => x"08",
          7726 => x"80",
          7727 => x"77",
          7728 => x"38",
          7729 => x"e4",
          7730 => x"0d",
          7731 => x"e4",
          7732 => x"b8",
          7733 => x"84",
          7734 => x"80",
          7735 => x"77",
          7736 => x"84",
          7737 => x"51",
          7738 => x"3f",
          7739 => x"e4",
          7740 => x"0d",
          7741 => x"f4",
          7742 => x"d4",
          7743 => x"0b",
          7744 => x"23",
          7745 => x"53",
          7746 => x"ff",
          7747 => x"b6",
          7748 => x"b8",
          7749 => x"76",
          7750 => x"0b",
          7751 => x"84",
          7752 => x"54",
          7753 => x"34",
          7754 => x"15",
          7755 => x"d4",
          7756 => x"86",
          7757 => x"0b",
          7758 => x"84",
          7759 => x"84",
          7760 => x"ff",
          7761 => x"80",
          7762 => x"ff",
          7763 => x"88",
          7764 => x"55",
          7765 => x"17",
          7766 => x"17",
          7767 => x"d0",
          7768 => x"10",
          7769 => x"d4",
          7770 => x"05",
          7771 => x"82",
          7772 => x"0b",
          7773 => x"77",
          7774 => x"2e",
          7775 => x"fe",
          7776 => x"3d",
          7777 => x"05",
          7778 => x"52",
          7779 => x"87",
          7780 => x"e0",
          7781 => x"71",
          7782 => x"0c",
          7783 => x"04",
          7784 => x"02",
          7785 => x"52",
          7786 => x"81",
          7787 => x"71",
          7788 => x"3f",
          7789 => x"08",
          7790 => x"53",
          7791 => x"72",
          7792 => x"13",
          7793 => x"e0",
          7794 => x"72",
          7795 => x"0c",
          7796 => x"04",
          7797 => x"7c",
          7798 => x"8c",
          7799 => x"33",
          7800 => x"59",
          7801 => x"74",
          7802 => x"84",
          7803 => x"33",
          7804 => x"06",
          7805 => x"73",
          7806 => x"58",
          7807 => x"c0",
          7808 => x"78",
          7809 => x"76",
          7810 => x"3f",
          7811 => x"08",
          7812 => x"55",
          7813 => x"a7",
          7814 => x"98",
          7815 => x"73",
          7816 => x"78",
          7817 => x"74",
          7818 => x"06",
          7819 => x"2e",
          7820 => x"54",
          7821 => x"84",
          7822 => x"8b",
          7823 => x"84",
          7824 => x"19",
          7825 => x"06",
          7826 => x"79",
          7827 => x"ac",
          7828 => x"f7",
          7829 => x"7e",
          7830 => x"05",
          7831 => x"5a",
          7832 => x"81",
          7833 => x"26",
          7834 => x"b8",
          7835 => x"54",
          7836 => x"54",
          7837 => x"bd",
          7838 => x"85",
          7839 => x"98",
          7840 => x"53",
          7841 => x"51",
          7842 => x"84",
          7843 => x"81",
          7844 => x"74",
          7845 => x"38",
          7846 => x"8c",
          7847 => x"e2",
          7848 => x"26",
          7849 => x"fc",
          7850 => x"54",
          7851 => x"83",
          7852 => x"73",
          7853 => x"b8",
          7854 => x"3d",
          7855 => x"80",
          7856 => x"70",
          7857 => x"5a",
          7858 => x"78",
          7859 => x"38",
          7860 => x"3d",
          7861 => x"84",
          7862 => x"33",
          7863 => x"9f",
          7864 => x"53",
          7865 => x"71",
          7866 => x"38",
          7867 => x"12",
          7868 => x"81",
          7869 => x"53",
          7870 => x"85",
          7871 => x"98",
          7872 => x"53",
          7873 => x"96",
          7874 => x"25",
          7875 => x"83",
          7876 => x"84",
          7877 => x"b8",
          7878 => x"3d",
          7879 => x"80",
          7880 => x"73",
          7881 => x"0c",
          7882 => x"04",
          7883 => x"0c",
          7884 => x"b8",
          7885 => x"3d",
          7886 => x"84",
          7887 => x"92",
          7888 => x"54",
          7889 => x"71",
          7890 => x"2a",
          7891 => x"51",
          7892 => x"8a",
          7893 => x"98",
          7894 => x"74",
          7895 => x"c0",
          7896 => x"51",
          7897 => x"81",
          7898 => x"c0",
          7899 => x"52",
          7900 => x"06",
          7901 => x"2e",
          7902 => x"71",
          7903 => x"54",
          7904 => x"ff",
          7905 => x"3d",
          7906 => x"80",
          7907 => x"33",
          7908 => x"57",
          7909 => x"09",
          7910 => x"38",
          7911 => x"75",
          7912 => x"87",
          7913 => x"80",
          7914 => x"33",
          7915 => x"3f",
          7916 => x"08",
          7917 => x"38",
          7918 => x"84",
          7919 => x"8c",
          7920 => x"81",
          7921 => x"08",
          7922 => x"70",
          7923 => x"33",
          7924 => x"ff",
          7925 => x"84",
          7926 => x"77",
          7927 => x"06",
          7928 => x"b8",
          7929 => x"19",
          7930 => x"08",
          7931 => x"08",
          7932 => x"08",
          7933 => x"08",
          7934 => x"5b",
          7935 => x"ff",
          7936 => x"18",
          7937 => x"82",
          7938 => x"06",
          7939 => x"81",
          7940 => x"53",
          7941 => x"18",
          7942 => x"b7",
          7943 => x"33",
          7944 => x"83",
          7945 => x"06",
          7946 => x"84",
          7947 => x"76",
          7948 => x"81",
          7949 => x"38",
          7950 => x"84",
          7951 => x"57",
          7952 => x"81",
          7953 => x"ff",
          7954 => x"f4",
          7955 => x"0b",
          7956 => x"34",
          7957 => x"84",
          7958 => x"80",
          7959 => x"80",
          7960 => x"19",
          7961 => x"0b",
          7962 => x"80",
          7963 => x"19",
          7964 => x"0b",
          7965 => x"34",
          7966 => x"84",
          7967 => x"80",
          7968 => x"9e",
          7969 => x"e1",
          7970 => x"19",
          7971 => x"08",
          7972 => x"a0",
          7973 => x"88",
          7974 => x"84",
          7975 => x"74",
          7976 => x"75",
          7977 => x"34",
          7978 => x"5b",
          7979 => x"19",
          7980 => x"08",
          7981 => x"a4",
          7982 => x"88",
          7983 => x"84",
          7984 => x"7a",
          7985 => x"75",
          7986 => x"34",
          7987 => x"55",
          7988 => x"19",
          7989 => x"08",
          7990 => x"b4",
          7991 => x"81",
          7992 => x"79",
          7993 => x"33",
          7994 => x"3f",
          7995 => x"34",
          7996 => x"52",
          7997 => x"51",
          7998 => x"84",
          7999 => x"80",
          8000 => x"38",
          8001 => x"f3",
          8002 => x"60",
          8003 => x"56",
          8004 => x"27",
          8005 => x"17",
          8006 => x"8c",
          8007 => x"77",
          8008 => x"0c",
          8009 => x"04",
          8010 => x"56",
          8011 => x"2e",
          8012 => x"74",
          8013 => x"a5",
          8014 => x"2e",
          8015 => x"dd",
          8016 => x"2a",
          8017 => x"2a",
          8018 => x"05",
          8019 => x"5b",
          8020 => x"79",
          8021 => x"83",
          8022 => x"7b",
          8023 => x"81",
          8024 => x"38",
          8025 => x"53",
          8026 => x"81",
          8027 => x"f8",
          8028 => x"b8",
          8029 => x"2e",
          8030 => x"59",
          8031 => x"b4",
          8032 => x"ff",
          8033 => x"83",
          8034 => x"b8",
          8035 => x"1c",
          8036 => x"a8",
          8037 => x"53",
          8038 => x"b4",
          8039 => x"2e",
          8040 => x"0b",
          8041 => x"71",
          8042 => x"74",
          8043 => x"81",
          8044 => x"38",
          8045 => x"53",
          8046 => x"81",
          8047 => x"f8",
          8048 => x"b8",
          8049 => x"2e",
          8050 => x"59",
          8051 => x"b4",
          8052 => x"fe",
          8053 => x"83",
          8054 => x"b8",
          8055 => x"88",
          8056 => x"78",
          8057 => x"84",
          8058 => x"59",
          8059 => x"fe",
          8060 => x"9f",
          8061 => x"b8",
          8062 => x"3d",
          8063 => x"88",
          8064 => x"08",
          8065 => x"17",
          8066 => x"b5",
          8067 => x"83",
          8068 => x"5c",
          8069 => x"7b",
          8070 => x"06",
          8071 => x"81",
          8072 => x"b8",
          8073 => x"17",
          8074 => x"a8",
          8075 => x"e4",
          8076 => x"85",
          8077 => x"81",
          8078 => x"18",
          8079 => x"df",
          8080 => x"83",
          8081 => x"05",
          8082 => x"11",
          8083 => x"71",
          8084 => x"84",
          8085 => x"57",
          8086 => x"0d",
          8087 => x"2e",
          8088 => x"fd",
          8089 => x"87",
          8090 => x"08",
          8091 => x"17",
          8092 => x"b5",
          8093 => x"83",
          8094 => x"5c",
          8095 => x"7b",
          8096 => x"06",
          8097 => x"81",
          8098 => x"b8",
          8099 => x"17",
          8100 => x"c0",
          8101 => x"e4",
          8102 => x"85",
          8103 => x"81",
          8104 => x"18",
          8105 => x"f7",
          8106 => x"2b",
          8107 => x"77",
          8108 => x"83",
          8109 => x"12",
          8110 => x"2b",
          8111 => x"07",
          8112 => x"70",
          8113 => x"2b",
          8114 => x"80",
          8115 => x"80",
          8116 => x"b8",
          8117 => x"5c",
          8118 => x"56",
          8119 => x"04",
          8120 => x"17",
          8121 => x"17",
          8122 => x"18",
          8123 => x"f6",
          8124 => x"5a",
          8125 => x"08",
          8126 => x"81",
          8127 => x"38",
          8128 => x"08",
          8129 => x"b4",
          8130 => x"18",
          8131 => x"b8",
          8132 => x"5e",
          8133 => x"08",
          8134 => x"38",
          8135 => x"55",
          8136 => x"09",
          8137 => x"f7",
          8138 => x"b4",
          8139 => x"18",
          8140 => x"7b",
          8141 => x"33",
          8142 => x"3f",
          8143 => x"df",
          8144 => x"b4",
          8145 => x"b8",
          8146 => x"81",
          8147 => x"5c",
          8148 => x"84",
          8149 => x"7b",
          8150 => x"06",
          8151 => x"84",
          8152 => x"83",
          8153 => x"17",
          8154 => x"08",
          8155 => x"a0",
          8156 => x"8b",
          8157 => x"33",
          8158 => x"2e",
          8159 => x"84",
          8160 => x"5b",
          8161 => x"81",
          8162 => x"08",
          8163 => x"70",
          8164 => x"33",
          8165 => x"bb",
          8166 => x"84",
          8167 => x"7b",
          8168 => x"06",
          8169 => x"84",
          8170 => x"83",
          8171 => x"17",
          8172 => x"08",
          8173 => x"e4",
          8174 => x"7d",
          8175 => x"27",
          8176 => x"82",
          8177 => x"74",
          8178 => x"81",
          8179 => x"38",
          8180 => x"17",
          8181 => x"08",
          8182 => x"52",
          8183 => x"51",
          8184 => x"7a",
          8185 => x"39",
          8186 => x"17",
          8187 => x"17",
          8188 => x"18",
          8189 => x"f4",
          8190 => x"5a",
          8191 => x"08",
          8192 => x"81",
          8193 => x"38",
          8194 => x"08",
          8195 => x"b4",
          8196 => x"18",
          8197 => x"b8",
          8198 => x"55",
          8199 => x"08",
          8200 => x"38",
          8201 => x"55",
          8202 => x"09",
          8203 => x"84",
          8204 => x"b4",
          8205 => x"18",
          8206 => x"7d",
          8207 => x"33",
          8208 => x"3f",
          8209 => x"ec",
          8210 => x"b4",
          8211 => x"18",
          8212 => x"7b",
          8213 => x"33",
          8214 => x"3f",
          8215 => x"81",
          8216 => x"bb",
          8217 => x"39",
          8218 => x"60",
          8219 => x"57",
          8220 => x"81",
          8221 => x"38",
          8222 => x"08",
          8223 => x"78",
          8224 => x"78",
          8225 => x"74",
          8226 => x"80",
          8227 => x"2e",
          8228 => x"77",
          8229 => x"0c",
          8230 => x"04",
          8231 => x"a8",
          8232 => x"58",
          8233 => x"1a",
          8234 => x"76",
          8235 => x"b6",
          8236 => x"33",
          8237 => x"7c",
          8238 => x"81",
          8239 => x"38",
          8240 => x"53",
          8241 => x"81",
          8242 => x"f2",
          8243 => x"b8",
          8244 => x"2e",
          8245 => x"58",
          8246 => x"b4",
          8247 => x"58",
          8248 => x"38",
          8249 => x"fe",
          8250 => x"7b",
          8251 => x"06",
          8252 => x"b8",
          8253 => x"88",
          8254 => x"b9",
          8255 => x"0b",
          8256 => x"77",
          8257 => x"0c",
          8258 => x"04",
          8259 => x"09",
          8260 => x"ff",
          8261 => x"2a",
          8262 => x"05",
          8263 => x"b4",
          8264 => x"5c",
          8265 => x"85",
          8266 => x"19",
          8267 => x"5d",
          8268 => x"09",
          8269 => x"bd",
          8270 => x"77",
          8271 => x"52",
          8272 => x"51",
          8273 => x"84",
          8274 => x"80",
          8275 => x"ff",
          8276 => x"77",
          8277 => x"79",
          8278 => x"b7",
          8279 => x"2b",
          8280 => x"79",
          8281 => x"83",
          8282 => x"98",
          8283 => x"06",
          8284 => x"06",
          8285 => x"5e",
          8286 => x"34",
          8287 => x"56",
          8288 => x"34",
          8289 => x"5a",
          8290 => x"34",
          8291 => x"5b",
          8292 => x"34",
          8293 => x"1a",
          8294 => x"39",
          8295 => x"16",
          8296 => x"a8",
          8297 => x"b4",
          8298 => x"59",
          8299 => x"2e",
          8300 => x"0b",
          8301 => x"71",
          8302 => x"74",
          8303 => x"81",
          8304 => x"38",
          8305 => x"53",
          8306 => x"81",
          8307 => x"f0",
          8308 => x"b8",
          8309 => x"2e",
          8310 => x"58",
          8311 => x"b4",
          8312 => x"58",
          8313 => x"38",
          8314 => x"06",
          8315 => x"81",
          8316 => x"06",
          8317 => x"7a",
          8318 => x"2e",
          8319 => x"84",
          8320 => x"06",
          8321 => x"06",
          8322 => x"5a",
          8323 => x"81",
          8324 => x"34",
          8325 => x"a8",
          8326 => x"56",
          8327 => x"1a",
          8328 => x"74",
          8329 => x"dd",
          8330 => x"74",
          8331 => x"70",
          8332 => x"33",
          8333 => x"9b",
          8334 => x"84",
          8335 => x"7f",
          8336 => x"06",
          8337 => x"84",
          8338 => x"83",
          8339 => x"19",
          8340 => x"1b",
          8341 => x"1b",
          8342 => x"e4",
          8343 => x"56",
          8344 => x"27",
          8345 => x"19",
          8346 => x"82",
          8347 => x"38",
          8348 => x"53",
          8349 => x"19",
          8350 => x"d8",
          8351 => x"e4",
          8352 => x"85",
          8353 => x"81",
          8354 => x"1a",
          8355 => x"83",
          8356 => x"ff",
          8357 => x"05",
          8358 => x"56",
          8359 => x"38",
          8360 => x"76",
          8361 => x"06",
          8362 => x"07",
          8363 => x"76",
          8364 => x"83",
          8365 => x"cb",
          8366 => x"76",
          8367 => x"70",
          8368 => x"33",
          8369 => x"8b",
          8370 => x"84",
          8371 => x"7c",
          8372 => x"06",
          8373 => x"84",
          8374 => x"83",
          8375 => x"19",
          8376 => x"1b",
          8377 => x"1b",
          8378 => x"e4",
          8379 => x"40",
          8380 => x"27",
          8381 => x"82",
          8382 => x"74",
          8383 => x"81",
          8384 => x"38",
          8385 => x"1e",
          8386 => x"81",
          8387 => x"ee",
          8388 => x"5a",
          8389 => x"81",
          8390 => x"b8",
          8391 => x"81",
          8392 => x"57",
          8393 => x"81",
          8394 => x"e4",
          8395 => x"09",
          8396 => x"ae",
          8397 => x"e4",
          8398 => x"34",
          8399 => x"70",
          8400 => x"31",
          8401 => x"84",
          8402 => x"5f",
          8403 => x"74",
          8404 => x"f0",
          8405 => x"33",
          8406 => x"2e",
          8407 => x"fc",
          8408 => x"54",
          8409 => x"76",
          8410 => x"33",
          8411 => x"3f",
          8412 => x"d0",
          8413 => x"76",
          8414 => x"70",
          8415 => x"33",
          8416 => x"cf",
          8417 => x"84",
          8418 => x"7c",
          8419 => x"06",
          8420 => x"84",
          8421 => x"83",
          8422 => x"19",
          8423 => x"1b",
          8424 => x"1b",
          8425 => x"e4",
          8426 => x"40",
          8427 => x"27",
          8428 => x"82",
          8429 => x"74",
          8430 => x"81",
          8431 => x"38",
          8432 => x"1e",
          8433 => x"81",
          8434 => x"ed",
          8435 => x"5a",
          8436 => x"81",
          8437 => x"53",
          8438 => x"19",
          8439 => x"f3",
          8440 => x"fd",
          8441 => x"76",
          8442 => x"06",
          8443 => x"83",
          8444 => x"59",
          8445 => x"b8",
          8446 => x"88",
          8447 => x"b9",
          8448 => x"fa",
          8449 => x"fd",
          8450 => x"76",
          8451 => x"fc",
          8452 => x"b8",
          8453 => x"33",
          8454 => x"8f",
          8455 => x"f0",
          8456 => x"42",
          8457 => x"58",
          8458 => x"7d",
          8459 => x"75",
          8460 => x"7d",
          8461 => x"79",
          8462 => x"7d",
          8463 => x"7a",
          8464 => x"fa",
          8465 => x"3d",
          8466 => x"71",
          8467 => x"5a",
          8468 => x"38",
          8469 => x"57",
          8470 => x"80",
          8471 => x"9c",
          8472 => x"80",
          8473 => x"19",
          8474 => x"54",
          8475 => x"80",
          8476 => x"7b",
          8477 => x"38",
          8478 => x"16",
          8479 => x"08",
          8480 => x"38",
          8481 => x"77",
          8482 => x"38",
          8483 => x"51",
          8484 => x"84",
          8485 => x"80",
          8486 => x"38",
          8487 => x"b8",
          8488 => x"2e",
          8489 => x"b8",
          8490 => x"70",
          8491 => x"07",
          8492 => x"7b",
          8493 => x"55",
          8494 => x"aa",
          8495 => x"2e",
          8496 => x"ff",
          8497 => x"55",
          8498 => x"e4",
          8499 => x"0d",
          8500 => x"ff",
          8501 => x"b8",
          8502 => x"ca",
          8503 => x"79",
          8504 => x"3f",
          8505 => x"84",
          8506 => x"27",
          8507 => x"b8",
          8508 => x"84",
          8509 => x"ff",
          8510 => x"9c",
          8511 => x"b8",
          8512 => x"c4",
          8513 => x"fe",
          8514 => x"1b",
          8515 => x"08",
          8516 => x"38",
          8517 => x"52",
          8518 => x"eb",
          8519 => x"84",
          8520 => x"81",
          8521 => x"38",
          8522 => x"08",
          8523 => x"70",
          8524 => x"25",
          8525 => x"84",
          8526 => x"54",
          8527 => x"55",
          8528 => x"38",
          8529 => x"08",
          8530 => x"38",
          8531 => x"54",
          8532 => x"fe",
          8533 => x"9c",
          8534 => x"fe",
          8535 => x"70",
          8536 => x"96",
          8537 => x"2e",
          8538 => x"ff",
          8539 => x"78",
          8540 => x"3f",
          8541 => x"08",
          8542 => x"08",
          8543 => x"b8",
          8544 => x"80",
          8545 => x"55",
          8546 => x"38",
          8547 => x"38",
          8548 => x"0c",
          8549 => x"fe",
          8550 => x"08",
          8551 => x"78",
          8552 => x"ff",
          8553 => x"0c",
          8554 => x"81",
          8555 => x"84",
          8556 => x"55",
          8557 => x"e4",
          8558 => x"0d",
          8559 => x"84",
          8560 => x"8c",
          8561 => x"84",
          8562 => x"58",
          8563 => x"73",
          8564 => x"b8",
          8565 => x"7a",
          8566 => x"f5",
          8567 => x"b8",
          8568 => x"ff",
          8569 => x"b8",
          8570 => x"b8",
          8571 => x"3d",
          8572 => x"56",
          8573 => x"ff",
          8574 => x"55",
          8575 => x"f8",
          8576 => x"7c",
          8577 => x"55",
          8578 => x"80",
          8579 => x"df",
          8580 => x"06",
          8581 => x"d7",
          8582 => x"19",
          8583 => x"08",
          8584 => x"df",
          8585 => x"56",
          8586 => x"80",
          8587 => x"85",
          8588 => x"0b",
          8589 => x"5a",
          8590 => x"27",
          8591 => x"17",
          8592 => x"0c",
          8593 => x"0c",
          8594 => x"53",
          8595 => x"80",
          8596 => x"73",
          8597 => x"98",
          8598 => x"83",
          8599 => x"b8",
          8600 => x"0c",
          8601 => x"84",
          8602 => x"8a",
          8603 => x"82",
          8604 => x"e4",
          8605 => x"0d",
          8606 => x"08",
          8607 => x"2e",
          8608 => x"8a",
          8609 => x"89",
          8610 => x"73",
          8611 => x"38",
          8612 => x"53",
          8613 => x"14",
          8614 => x"59",
          8615 => x"8d",
          8616 => x"22",
          8617 => x"b0",
          8618 => x"5a",
          8619 => x"19",
          8620 => x"39",
          8621 => x"51",
          8622 => x"84",
          8623 => x"55",
          8624 => x"08",
          8625 => x"38",
          8626 => x"b8",
          8627 => x"ff",
          8628 => x"17",
          8629 => x"b8",
          8630 => x"27",
          8631 => x"73",
          8632 => x"73",
          8633 => x"38",
          8634 => x"81",
          8635 => x"e4",
          8636 => x"0d",
          8637 => x"0d",
          8638 => x"90",
          8639 => x"05",
          8640 => x"f0",
          8641 => x"27",
          8642 => x"0b",
          8643 => x"98",
          8644 => x"84",
          8645 => x"2e",
          8646 => x"83",
          8647 => x"7a",
          8648 => x"15",
          8649 => x"57",
          8650 => x"38",
          8651 => x"88",
          8652 => x"55",
          8653 => x"81",
          8654 => x"98",
          8655 => x"90",
          8656 => x"1b",
          8657 => x"18",
          8658 => x"75",
          8659 => x"0c",
          8660 => x"04",
          8661 => x"0c",
          8662 => x"ff",
          8663 => x"2a",
          8664 => x"da",
          8665 => x"76",
          8666 => x"3f",
          8667 => x"08",
          8668 => x"81",
          8669 => x"e4",
          8670 => x"38",
          8671 => x"b8",
          8672 => x"2e",
          8673 => x"19",
          8674 => x"e4",
          8675 => x"91",
          8676 => x"2e",
          8677 => x"94",
          8678 => x"76",
          8679 => x"3f",
          8680 => x"08",
          8681 => x"84",
          8682 => x"80",
          8683 => x"38",
          8684 => x"b8",
          8685 => x"2e",
          8686 => x"81",
          8687 => x"e4",
          8688 => x"ff",
          8689 => x"b8",
          8690 => x"1a",
          8691 => x"7d",
          8692 => x"fe",
          8693 => x"08",
          8694 => x"56",
          8695 => x"78",
          8696 => x"8a",
          8697 => x"71",
          8698 => x"08",
          8699 => x"7b",
          8700 => x"b8",
          8701 => x"80",
          8702 => x"80",
          8703 => x"05",
          8704 => x"15",
          8705 => x"38",
          8706 => x"19",
          8707 => x"75",
          8708 => x"38",
          8709 => x"1c",
          8710 => x"81",
          8711 => x"e4",
          8712 => x"b8",
          8713 => x"e7",
          8714 => x"56",
          8715 => x"98",
          8716 => x"0b",
          8717 => x"0c",
          8718 => x"04",
          8719 => x"19",
          8720 => x"19",
          8721 => x"1a",
          8722 => x"e4",
          8723 => x"b8",
          8724 => x"f3",
          8725 => x"e4",
          8726 => x"34",
          8727 => x"a8",
          8728 => x"55",
          8729 => x"08",
          8730 => x"38",
          8731 => x"5c",
          8732 => x"09",
          8733 => x"db",
          8734 => x"b4",
          8735 => x"1a",
          8736 => x"75",
          8737 => x"33",
          8738 => x"3f",
          8739 => x"8a",
          8740 => x"74",
          8741 => x"06",
          8742 => x"2e",
          8743 => x"a7",
          8744 => x"18",
          8745 => x"9c",
          8746 => x"05",
          8747 => x"58",
          8748 => x"fd",
          8749 => x"19",
          8750 => x"29",
          8751 => x"05",
          8752 => x"5c",
          8753 => x"81",
          8754 => x"e4",
          8755 => x"0d",
          8756 => x"0d",
          8757 => x"5c",
          8758 => x"5a",
          8759 => x"70",
          8760 => x"58",
          8761 => x"80",
          8762 => x"38",
          8763 => x"75",
          8764 => x"b4",
          8765 => x"2e",
          8766 => x"83",
          8767 => x"58",
          8768 => x"2e",
          8769 => x"81",
          8770 => x"54",
          8771 => x"19",
          8772 => x"33",
          8773 => x"3f",
          8774 => x"08",
          8775 => x"38",
          8776 => x"57",
          8777 => x"0c",
          8778 => x"82",
          8779 => x"1c",
          8780 => x"58",
          8781 => x"2e",
          8782 => x"8b",
          8783 => x"06",
          8784 => x"06",
          8785 => x"86",
          8786 => x"81",
          8787 => x"30",
          8788 => x"70",
          8789 => x"25",
          8790 => x"07",
          8791 => x"57",
          8792 => x"38",
          8793 => x"06",
          8794 => x"88",
          8795 => x"38",
          8796 => x"81",
          8797 => x"ff",
          8798 => x"7b",
          8799 => x"3f",
          8800 => x"08",
          8801 => x"e4",
          8802 => x"38",
          8803 => x"56",
          8804 => x"38",
          8805 => x"e4",
          8806 => x"0d",
          8807 => x"b4",
          8808 => x"7e",
          8809 => x"33",
          8810 => x"3f",
          8811 => x"b8",
          8812 => x"2e",
          8813 => x"fe",
          8814 => x"b8",
          8815 => x"1a",
          8816 => x"08",
          8817 => x"31",
          8818 => x"08",
          8819 => x"a0",
          8820 => x"fe",
          8821 => x"19",
          8822 => x"82",
          8823 => x"06",
          8824 => x"81",
          8825 => x"08",
          8826 => x"05",
          8827 => x"81",
          8828 => x"e0",
          8829 => x"57",
          8830 => x"79",
          8831 => x"81",
          8832 => x"38",
          8833 => x"81",
          8834 => x"80",
          8835 => x"8d",
          8836 => x"81",
          8837 => x"90",
          8838 => x"ac",
          8839 => x"5e",
          8840 => x"2e",
          8841 => x"ff",
          8842 => x"fe",
          8843 => x"56",
          8844 => x"09",
          8845 => x"be",
          8846 => x"84",
          8847 => x"98",
          8848 => x"84",
          8849 => x"94",
          8850 => x"77",
          8851 => x"39",
          8852 => x"57",
          8853 => x"09",
          8854 => x"38",
          8855 => x"9b",
          8856 => x"1a",
          8857 => x"2b",
          8858 => x"41",
          8859 => x"38",
          8860 => x"81",
          8861 => x"29",
          8862 => x"5a",
          8863 => x"5b",
          8864 => x"17",
          8865 => x"81",
          8866 => x"33",
          8867 => x"07",
          8868 => x"7a",
          8869 => x"c5",
          8870 => x"fe",
          8871 => x"38",
          8872 => x"05",
          8873 => x"75",
          8874 => x"1a",
          8875 => x"57",
          8876 => x"cc",
          8877 => x"70",
          8878 => x"06",
          8879 => x"80",
          8880 => x"79",
          8881 => x"fe",
          8882 => x"10",
          8883 => x"80",
          8884 => x"1d",
          8885 => x"06",
          8886 => x"9d",
          8887 => x"ff",
          8888 => x"38",
          8889 => x"fe",
          8890 => x"a8",
          8891 => x"8b",
          8892 => x"2a",
          8893 => x"29",
          8894 => x"81",
          8895 => x"40",
          8896 => x"81",
          8897 => x"19",
          8898 => x"76",
          8899 => x"7e",
          8900 => x"38",
          8901 => x"1d",
          8902 => x"b8",
          8903 => x"3d",
          8904 => x"3d",
          8905 => x"08",
          8906 => x"52",
          8907 => x"cf",
          8908 => x"e4",
          8909 => x"b8",
          8910 => x"80",
          8911 => x"70",
          8912 => x"0b",
          8913 => x"b8",
          8914 => x"1c",
          8915 => x"58",
          8916 => x"76",
          8917 => x"38",
          8918 => x"78",
          8919 => x"78",
          8920 => x"06",
          8921 => x"81",
          8922 => x"b8",
          8923 => x"1b",
          8924 => x"e0",
          8925 => x"e4",
          8926 => x"85",
          8927 => x"81",
          8928 => x"1c",
          8929 => x"76",
          8930 => x"9c",
          8931 => x"33",
          8932 => x"80",
          8933 => x"38",
          8934 => x"bf",
          8935 => x"ff",
          8936 => x"77",
          8937 => x"76",
          8938 => x"80",
          8939 => x"83",
          8940 => x"55",
          8941 => x"81",
          8942 => x"80",
          8943 => x"8f",
          8944 => x"38",
          8945 => x"78",
          8946 => x"8b",
          8947 => x"2a",
          8948 => x"29",
          8949 => x"81",
          8950 => x"57",
          8951 => x"81",
          8952 => x"19",
          8953 => x"76",
          8954 => x"7f",
          8955 => x"38",
          8956 => x"81",
          8957 => x"a7",
          8958 => x"a0",
          8959 => x"78",
          8960 => x"5a",
          8961 => x"81",
          8962 => x"71",
          8963 => x"1a",
          8964 => x"40",
          8965 => x"81",
          8966 => x"80",
          8967 => x"81",
          8968 => x"0b",
          8969 => x"80",
          8970 => x"f5",
          8971 => x"b8",
          8972 => x"84",
          8973 => x"80",
          8974 => x"38",
          8975 => x"e4",
          8976 => x"0d",
          8977 => x"b4",
          8978 => x"7d",
          8979 => x"33",
          8980 => x"3f",
          8981 => x"b8",
          8982 => x"2e",
          8983 => x"fe",
          8984 => x"b8",
          8985 => x"1c",
          8986 => x"08",
          8987 => x"31",
          8988 => x"08",
          8989 => x"a0",
          8990 => x"fd",
          8991 => x"1b",
          8992 => x"82",
          8993 => x"06",
          8994 => x"81",
          8995 => x"08",
          8996 => x"05",
          8997 => x"81",
          8998 => x"db",
          8999 => x"57",
          9000 => x"77",
          9001 => x"39",
          9002 => x"70",
          9003 => x"06",
          9004 => x"fe",
          9005 => x"86",
          9006 => x"5a",
          9007 => x"93",
          9008 => x"33",
          9009 => x"06",
          9010 => x"08",
          9011 => x"0c",
          9012 => x"76",
          9013 => x"38",
          9014 => x"74",
          9015 => x"7b",
          9016 => x"3f",
          9017 => x"08",
          9018 => x"e4",
          9019 => x"fc",
          9020 => x"c8",
          9021 => x"2e",
          9022 => x"81",
          9023 => x"0b",
          9024 => x"fe",
          9025 => x"19",
          9026 => x"77",
          9027 => x"06",
          9028 => x"1b",
          9029 => x"33",
          9030 => x"71",
          9031 => x"59",
          9032 => x"ff",
          9033 => x"33",
          9034 => x"8d",
          9035 => x"5b",
          9036 => x"59",
          9037 => x"e4",
          9038 => x"05",
          9039 => x"71",
          9040 => x"2b",
          9041 => x"57",
          9042 => x"80",
          9043 => x"81",
          9044 => x"84",
          9045 => x"81",
          9046 => x"84",
          9047 => x"7a",
          9048 => x"70",
          9049 => x"81",
          9050 => x"81",
          9051 => x"75",
          9052 => x"08",
          9053 => x"06",
          9054 => x"76",
          9055 => x"58",
          9056 => x"ff",
          9057 => x"33",
          9058 => x"81",
          9059 => x"75",
          9060 => x"38",
          9061 => x"8d",
          9062 => x"60",
          9063 => x"41",
          9064 => x"b4",
          9065 => x"70",
          9066 => x"5e",
          9067 => x"39",
          9068 => x"b8",
          9069 => x"3d",
          9070 => x"83",
          9071 => x"ff",
          9072 => x"ff",
          9073 => x"39",
          9074 => x"68",
          9075 => x"ab",
          9076 => x"a0",
          9077 => x"5d",
          9078 => x"74",
          9079 => x"74",
          9080 => x"70",
          9081 => x"5d",
          9082 => x"8e",
          9083 => x"70",
          9084 => x"22",
          9085 => x"74",
          9086 => x"3d",
          9087 => x"40",
          9088 => x"58",
          9089 => x"70",
          9090 => x"33",
          9091 => x"05",
          9092 => x"15",
          9093 => x"38",
          9094 => x"05",
          9095 => x"06",
          9096 => x"80",
          9097 => x"38",
          9098 => x"ab",
          9099 => x"0b",
          9100 => x"5b",
          9101 => x"7b",
          9102 => x"7a",
          9103 => x"55",
          9104 => x"05",
          9105 => x"70",
          9106 => x"34",
          9107 => x"74",
          9108 => x"7b",
          9109 => x"38",
          9110 => x"56",
          9111 => x"2e",
          9112 => x"82",
          9113 => x"8f",
          9114 => x"06",
          9115 => x"76",
          9116 => x"83",
          9117 => x"72",
          9118 => x"06",
          9119 => x"57",
          9120 => x"87",
          9121 => x"a0",
          9122 => x"ff",
          9123 => x"80",
          9124 => x"78",
          9125 => x"ca",
          9126 => x"84",
          9127 => x"05",
          9128 => x"b0",
          9129 => x"55",
          9130 => x"84",
          9131 => x"55",
          9132 => x"ff",
          9133 => x"78",
          9134 => x"59",
          9135 => x"38",
          9136 => x"80",
          9137 => x"76",
          9138 => x"80",
          9139 => x"38",
          9140 => x"74",
          9141 => x"38",
          9142 => x"75",
          9143 => x"a2",
          9144 => x"70",
          9145 => x"74",
          9146 => x"81",
          9147 => x"81",
          9148 => x"55",
          9149 => x"8e",
          9150 => x"78",
          9151 => x"81",
          9152 => x"57",
          9153 => x"77",
          9154 => x"27",
          9155 => x"7d",
          9156 => x"3f",
          9157 => x"08",
          9158 => x"1b",
          9159 => x"7b",
          9160 => x"38",
          9161 => x"80",
          9162 => x"e7",
          9163 => x"e4",
          9164 => x"b8",
          9165 => x"2e",
          9166 => x"82",
          9167 => x"80",
          9168 => x"ab",
          9169 => x"08",
          9170 => x"80",
          9171 => x"57",
          9172 => x"2a",
          9173 => x"81",
          9174 => x"2e",
          9175 => x"52",
          9176 => x"fe",
          9177 => x"84",
          9178 => x"1b",
          9179 => x"7d",
          9180 => x"3f",
          9181 => x"08",
          9182 => x"e4",
          9183 => x"38",
          9184 => x"08",
          9185 => x"59",
          9186 => x"56",
          9187 => x"18",
          9188 => x"85",
          9189 => x"18",
          9190 => x"77",
          9191 => x"06",
          9192 => x"81",
          9193 => x"b8",
          9194 => x"18",
          9195 => x"a4",
          9196 => x"e4",
          9197 => x"85",
          9198 => x"81",
          9199 => x"19",
          9200 => x"76",
          9201 => x"1e",
          9202 => x"56",
          9203 => x"e5",
          9204 => x"38",
          9205 => x"80",
          9206 => x"56",
          9207 => x"2e",
          9208 => x"81",
          9209 => x"7b",
          9210 => x"38",
          9211 => x"51",
          9212 => x"84",
          9213 => x"56",
          9214 => x"08",
          9215 => x"88",
          9216 => x"75",
          9217 => x"89",
          9218 => x"75",
          9219 => x"ff",
          9220 => x"81",
          9221 => x"1e",
          9222 => x"1c",
          9223 => x"af",
          9224 => x"33",
          9225 => x"7f",
          9226 => x"81",
          9227 => x"b8",
          9228 => x"1c",
          9229 => x"9c",
          9230 => x"e4",
          9231 => x"85",
          9232 => x"81",
          9233 => x"1d",
          9234 => x"75",
          9235 => x"a0",
          9236 => x"08",
          9237 => x"76",
          9238 => x"58",
          9239 => x"55",
          9240 => x"8b",
          9241 => x"08",
          9242 => x"55",
          9243 => x"05",
          9244 => x"70",
          9245 => x"34",
          9246 => x"74",
          9247 => x"1e",
          9248 => x"33",
          9249 => x"5a",
          9250 => x"34",
          9251 => x"1d",
          9252 => x"75",
          9253 => x"0c",
          9254 => x"04",
          9255 => x"70",
          9256 => x"07",
          9257 => x"74",
          9258 => x"74",
          9259 => x"7d",
          9260 => x"3f",
          9261 => x"08",
          9262 => x"e4",
          9263 => x"fd",
          9264 => x"bd",
          9265 => x"b4",
          9266 => x"7c",
          9267 => x"33",
          9268 => x"3f",
          9269 => x"08",
          9270 => x"81",
          9271 => x"38",
          9272 => x"08",
          9273 => x"b4",
          9274 => x"19",
          9275 => x"74",
          9276 => x"27",
          9277 => x"18",
          9278 => x"82",
          9279 => x"38",
          9280 => x"08",
          9281 => x"39",
          9282 => x"90",
          9283 => x"31",
          9284 => x"51",
          9285 => x"84",
          9286 => x"58",
          9287 => x"08",
          9288 => x"79",
          9289 => x"08",
          9290 => x"57",
          9291 => x"75",
          9292 => x"05",
          9293 => x"05",
          9294 => x"76",
          9295 => x"ff",
          9296 => x"59",
          9297 => x"e4",
          9298 => x"ff",
          9299 => x"43",
          9300 => x"08",
          9301 => x"b4",
          9302 => x"2e",
          9303 => x"1c",
          9304 => x"76",
          9305 => x"06",
          9306 => x"81",
          9307 => x"b8",
          9308 => x"1c",
          9309 => x"dc",
          9310 => x"e4",
          9311 => x"85",
          9312 => x"81",
          9313 => x"1d",
          9314 => x"75",
          9315 => x"8c",
          9316 => x"1f",
          9317 => x"ff",
          9318 => x"5f",
          9319 => x"34",
          9320 => x"1c",
          9321 => x"1c",
          9322 => x"1c",
          9323 => x"1c",
          9324 => x"29",
          9325 => x"77",
          9326 => x"76",
          9327 => x"2e",
          9328 => x"10",
          9329 => x"81",
          9330 => x"56",
          9331 => x"18",
          9332 => x"55",
          9333 => x"81",
          9334 => x"76",
          9335 => x"75",
          9336 => x"85",
          9337 => x"ff",
          9338 => x"58",
          9339 => x"cb",
          9340 => x"ff",
          9341 => x"b3",
          9342 => x"1f",
          9343 => x"58",
          9344 => x"81",
          9345 => x"7b",
          9346 => x"83",
          9347 => x"52",
          9348 => x"e1",
          9349 => x"e4",
          9350 => x"b8",
          9351 => x"f1",
          9352 => x"05",
          9353 => x"a9",
          9354 => x"39",
          9355 => x"1c",
          9356 => x"1c",
          9357 => x"1d",
          9358 => x"d0",
          9359 => x"56",
          9360 => x"08",
          9361 => x"84",
          9362 => x"83",
          9363 => x"1c",
          9364 => x"08",
          9365 => x"e4",
          9366 => x"60",
          9367 => x"27",
          9368 => x"82",
          9369 => x"61",
          9370 => x"81",
          9371 => x"38",
          9372 => x"1c",
          9373 => x"08",
          9374 => x"52",
          9375 => x"51",
          9376 => x"77",
          9377 => x"39",
          9378 => x"08",
          9379 => x"43",
          9380 => x"e5",
          9381 => x"06",
          9382 => x"fb",
          9383 => x"70",
          9384 => x"80",
          9385 => x"38",
          9386 => x"7c",
          9387 => x"5d",
          9388 => x"81",
          9389 => x"08",
          9390 => x"81",
          9391 => x"cf",
          9392 => x"b8",
          9393 => x"2e",
          9394 => x"bc",
          9395 => x"e4",
          9396 => x"34",
          9397 => x"a8",
          9398 => x"55",
          9399 => x"08",
          9400 => x"82",
          9401 => x"7e",
          9402 => x"38",
          9403 => x"08",
          9404 => x"39",
          9405 => x"41",
          9406 => x"2e",
          9407 => x"fc",
          9408 => x"1a",
          9409 => x"39",
          9410 => x"56",
          9411 => x"fc",
          9412 => x"fd",
          9413 => x"b4",
          9414 => x"1d",
          9415 => x"61",
          9416 => x"33",
          9417 => x"3f",
          9418 => x"81",
          9419 => x"08",
          9420 => x"05",
          9421 => x"81",
          9422 => x"ce",
          9423 => x"e3",
          9424 => x"0d",
          9425 => x"08",
          9426 => x"80",
          9427 => x"34",
          9428 => x"80",
          9429 => x"38",
          9430 => x"ff",
          9431 => x"38",
          9432 => x"60",
          9433 => x"70",
          9434 => x"5b",
          9435 => x"78",
          9436 => x"77",
          9437 => x"70",
          9438 => x"5b",
          9439 => x"82",
          9440 => x"d0",
          9441 => x"83",
          9442 => x"58",
          9443 => x"ff",
          9444 => x"38",
          9445 => x"76",
          9446 => x"5d",
          9447 => x"79",
          9448 => x"30",
          9449 => x"70",
          9450 => x"5a",
          9451 => x"18",
          9452 => x"80",
          9453 => x"34",
          9454 => x"1f",
          9455 => x"9c",
          9456 => x"70",
          9457 => x"58",
          9458 => x"a0",
          9459 => x"74",
          9460 => x"bc",
          9461 => x"32",
          9462 => x"72",
          9463 => x"55",
          9464 => x"8b",
          9465 => x"72",
          9466 => x"38",
          9467 => x"81",
          9468 => x"81",
          9469 => x"77",
          9470 => x"59",
          9471 => x"58",
          9472 => x"ff",
          9473 => x"18",
          9474 => x"80",
          9475 => x"34",
          9476 => x"53",
          9477 => x"77",
          9478 => x"bf",
          9479 => x"34",
          9480 => x"17",
          9481 => x"80",
          9482 => x"34",
          9483 => x"8c",
          9484 => x"53",
          9485 => x"73",
          9486 => x"9c",
          9487 => x"8b",
          9488 => x"1e",
          9489 => x"08",
          9490 => x"11",
          9491 => x"33",
          9492 => x"71",
          9493 => x"81",
          9494 => x"72",
          9495 => x"75",
          9496 => x"64",
          9497 => x"16",
          9498 => x"33",
          9499 => x"07",
          9500 => x"40",
          9501 => x"55",
          9502 => x"23",
          9503 => x"98",
          9504 => x"88",
          9505 => x"54",
          9506 => x"23",
          9507 => x"04",
          9508 => x"fe",
          9509 => x"1d",
          9510 => x"ff",
          9511 => x"5b",
          9512 => x"52",
          9513 => x"74",
          9514 => x"91",
          9515 => x"b8",
          9516 => x"ff",
          9517 => x"81",
          9518 => x"ad",
          9519 => x"27",
          9520 => x"74",
          9521 => x"73",
          9522 => x"97",
          9523 => x"78",
          9524 => x"0b",
          9525 => x"56",
          9526 => x"75",
          9527 => x"5c",
          9528 => x"fd",
          9529 => x"ba",
          9530 => x"76",
          9531 => x"07",
          9532 => x"80",
          9533 => x"55",
          9534 => x"f9",
          9535 => x"34",
          9536 => x"58",
          9537 => x"1f",
          9538 => x"cd",
          9539 => x"89",
          9540 => x"57",
          9541 => x"2e",
          9542 => x"7c",
          9543 => x"57",
          9544 => x"14",
          9545 => x"11",
          9546 => x"99",
          9547 => x"9c",
          9548 => x"11",
          9549 => x"88",
          9550 => x"38",
          9551 => x"53",
          9552 => x"5e",
          9553 => x"8a",
          9554 => x"70",
          9555 => x"06",
          9556 => x"78",
          9557 => x"5a",
          9558 => x"81",
          9559 => x"71",
          9560 => x"5e",
          9561 => x"56",
          9562 => x"38",
          9563 => x"72",
          9564 => x"cc",
          9565 => x"30",
          9566 => x"70",
          9567 => x"53",
          9568 => x"fc",
          9569 => x"3d",
          9570 => x"08",
          9571 => x"5c",
          9572 => x"33",
          9573 => x"74",
          9574 => x"38",
          9575 => x"80",
          9576 => x"df",
          9577 => x"2e",
          9578 => x"98",
          9579 => x"1d",
          9580 => x"96",
          9581 => x"41",
          9582 => x"75",
          9583 => x"38",
          9584 => x"16",
          9585 => x"57",
          9586 => x"81",
          9587 => x"55",
          9588 => x"df",
          9589 => x"0c",
          9590 => x"81",
          9591 => x"ff",
          9592 => x"8b",
          9593 => x"18",
          9594 => x"23",
          9595 => x"73",
          9596 => x"06",
          9597 => x"70",
          9598 => x"27",
          9599 => x"07",
          9600 => x"55",
          9601 => x"38",
          9602 => x"2e",
          9603 => x"74",
          9604 => x"b2",
          9605 => x"80",
          9606 => x"80",
          9607 => x"ff",
          9608 => x"56",
          9609 => x"81",
          9610 => x"75",
          9611 => x"81",
          9612 => x"70",
          9613 => x"56",
          9614 => x"ee",
          9615 => x"ff",
          9616 => x"81",
          9617 => x"81",
          9618 => x"fd",
          9619 => x"18",
          9620 => x"23",
          9621 => x"70",
          9622 => x"52",
          9623 => x"57",
          9624 => x"fe",
          9625 => x"cb",
          9626 => x"80",
          9627 => x"30",
          9628 => x"73",
          9629 => x"58",
          9630 => x"2e",
          9631 => x"14",
          9632 => x"80",
          9633 => x"55",
          9634 => x"dd",
          9635 => x"dc",
          9636 => x"70",
          9637 => x"07",
          9638 => x"72",
          9639 => x"88",
          9640 => x"33",
          9641 => x"3d",
          9642 => x"74",
          9643 => x"90",
          9644 => x"83",
          9645 => x"51",
          9646 => x"3f",
          9647 => x"08",
          9648 => x"06",
          9649 => x"8d",
          9650 => x"73",
          9651 => x"0c",
          9652 => x"04",
          9653 => x"33",
          9654 => x"06",
          9655 => x"80",
          9656 => x"38",
          9657 => x"80",
          9658 => x"34",
          9659 => x"51",
          9660 => x"84",
          9661 => x"84",
          9662 => x"93",
          9663 => x"81",
          9664 => x"32",
          9665 => x"80",
          9666 => x"41",
          9667 => x"7d",
          9668 => x"38",
          9669 => x"80",
          9670 => x"55",
          9671 => x"af",
          9672 => x"72",
          9673 => x"70",
          9674 => x"25",
          9675 => x"54",
          9676 => x"38",
          9677 => x"9f",
          9678 => x"2b",
          9679 => x"2e",
          9680 => x"76",
          9681 => x"d1",
          9682 => x"59",
          9683 => x"a7",
          9684 => x"78",
          9685 => x"70",
          9686 => x"32",
          9687 => x"9f",
          9688 => x"56",
          9689 => x"7c",
          9690 => x"38",
          9691 => x"ff",
          9692 => x"dd",
          9693 => x"77",
          9694 => x"76",
          9695 => x"2e",
          9696 => x"80",
          9697 => x"83",
          9698 => x"72",
          9699 => x"56",
          9700 => x"82",
          9701 => x"83",
          9702 => x"53",
          9703 => x"82",
          9704 => x"80",
          9705 => x"77",
          9706 => x"70",
          9707 => x"78",
          9708 => x"38",
          9709 => x"fe",
          9710 => x"17",
          9711 => x"2e",
          9712 => x"14",
          9713 => x"54",
          9714 => x"09",
          9715 => x"38",
          9716 => x"1d",
          9717 => x"74",
          9718 => x"56",
          9719 => x"53",
          9720 => x"72",
          9721 => x"88",
          9722 => x"22",
          9723 => x"57",
          9724 => x"80",
          9725 => x"38",
          9726 => x"83",
          9727 => x"ae",
          9728 => x"70",
          9729 => x"5a",
          9730 => x"2e",
          9731 => x"72",
          9732 => x"72",
          9733 => x"26",
          9734 => x"59",
          9735 => x"70",
          9736 => x"07",
          9737 => x"7c",
          9738 => x"54",
          9739 => x"2e",
          9740 => x"7c",
          9741 => x"83",
          9742 => x"2e",
          9743 => x"83",
          9744 => x"77",
          9745 => x"76",
          9746 => x"8b",
          9747 => x"81",
          9748 => x"18",
          9749 => x"77",
          9750 => x"81",
          9751 => x"53",
          9752 => x"38",
          9753 => x"57",
          9754 => x"2e",
          9755 => x"7c",
          9756 => x"e3",
          9757 => x"06",
          9758 => x"2e",
          9759 => x"7d",
          9760 => x"74",
          9761 => x"e3",
          9762 => x"2a",
          9763 => x"75",
          9764 => x"81",
          9765 => x"80",
          9766 => x"79",
          9767 => x"7d",
          9768 => x"06",
          9769 => x"2e",
          9770 => x"88",
          9771 => x"ab",
          9772 => x"51",
          9773 => x"84",
          9774 => x"ab",
          9775 => x"54",
          9776 => x"08",
          9777 => x"ac",
          9778 => x"e4",
          9779 => x"09",
          9780 => x"f7",
          9781 => x"2a",
          9782 => x"79",
          9783 => x"f0",
          9784 => x"2a",
          9785 => x"78",
          9786 => x"7b",
          9787 => x"56",
          9788 => x"16",
          9789 => x"57",
          9790 => x"81",
          9791 => x"79",
          9792 => x"40",
          9793 => x"7c",
          9794 => x"38",
          9795 => x"fd",
          9796 => x"83",
          9797 => x"8a",
          9798 => x"22",
          9799 => x"2e",
          9800 => x"fc",
          9801 => x"22",
          9802 => x"2e",
          9803 => x"fc",
          9804 => x"10",
          9805 => x"7b",
          9806 => x"a0",
          9807 => x"ae",
          9808 => x"26",
          9809 => x"54",
          9810 => x"81",
          9811 => x"81",
          9812 => x"73",
          9813 => x"79",
          9814 => x"77",
          9815 => x"7b",
          9816 => x"3f",
          9817 => x"08",
          9818 => x"56",
          9819 => x"e4",
          9820 => x"38",
          9821 => x"81",
          9822 => x"fa",
          9823 => x"1c",
          9824 => x"2a",
          9825 => x"5d",
          9826 => x"83",
          9827 => x"1c",
          9828 => x"06",
          9829 => x"d3",
          9830 => x"d2",
          9831 => x"88",
          9832 => x"33",
          9833 => x"54",
          9834 => x"82",
          9835 => x"88",
          9836 => x"08",
          9837 => x"fe",
          9838 => x"22",
          9839 => x"2e",
          9840 => x"76",
          9841 => x"fb",
          9842 => x"ab",
          9843 => x"07",
          9844 => x"5a",
          9845 => x"7d",
          9846 => x"fc",
          9847 => x"06",
          9848 => x"8c",
          9849 => x"06",
          9850 => x"79",
          9851 => x"fd",
          9852 => x"0b",
          9853 => x"7c",
          9854 => x"81",
          9855 => x"38",
          9856 => x"80",
          9857 => x"34",
          9858 => x"b8",
          9859 => x"3d",
          9860 => x"80",
          9861 => x"38",
          9862 => x"27",
          9863 => x"ff",
          9864 => x"7b",
          9865 => x"38",
          9866 => x"7d",
          9867 => x"5c",
          9868 => x"39",
          9869 => x"5a",
          9870 => x"74",
          9871 => x"f6",
          9872 => x"e4",
          9873 => x"ff",
          9874 => x"2a",
          9875 => x"55",
          9876 => x"c4",
          9877 => x"ff",
          9878 => x"f4",
          9879 => x"54",
          9880 => x"26",
          9881 => x"74",
          9882 => x"85",
          9883 => x"8c",
          9884 => x"8c",
          9885 => x"ff",
          9886 => x"59",
          9887 => x"80",
          9888 => x"75",
          9889 => x"81",
          9890 => x"70",
          9891 => x"56",
          9892 => x"ee",
          9893 => x"ff",
          9894 => x"80",
          9895 => x"bf",
          9896 => x"99",
          9897 => x"7d",
          9898 => x"81",
          9899 => x"53",
          9900 => x"59",
          9901 => x"93",
          9902 => x"07",
          9903 => x"06",
          9904 => x"83",
          9905 => x"58",
          9906 => x"7b",
          9907 => x"59",
          9908 => x"81",
          9909 => x"16",
          9910 => x"39",
          9911 => x"b3",
          9912 => x"8c",
          9913 => x"ff",
          9914 => x"78",
          9915 => x"ae",
          9916 => x"7a",
          9917 => x"1d",
          9918 => x"5b",
          9919 => x"34",
          9920 => x"d2",
          9921 => x"14",
          9922 => x"15",
          9923 => x"2b",
          9924 => x"07",
          9925 => x"1f",
          9926 => x"fd",
          9927 => x"1b",
          9928 => x"88",
          9929 => x"72",
          9930 => x"1b",
          9931 => x"05",
          9932 => x"79",
          9933 => x"5b",
          9934 => x"79",
          9935 => x"1d",
          9936 => x"76",
          9937 => x"09",
          9938 => x"a3",
          9939 => x"39",
          9940 => x"81",
          9941 => x"f6",
          9942 => x"0b",
          9943 => x"0c",
          9944 => x"04",
          9945 => x"67",
          9946 => x"05",
          9947 => x"33",
          9948 => x"80",
          9949 => x"7e",
          9950 => x"5b",
          9951 => x"2e",
          9952 => x"79",
          9953 => x"5b",
          9954 => x"26",
          9955 => x"ba",
          9956 => x"38",
          9957 => x"75",
          9958 => x"c7",
          9959 => x"c0",
          9960 => x"76",
          9961 => x"38",
          9962 => x"84",
          9963 => x"70",
          9964 => x"8c",
          9965 => x"2e",
          9966 => x"76",
          9967 => x"81",
          9968 => x"33",
          9969 => x"80",
          9970 => x"81",
          9971 => x"ff",
          9972 => x"84",
          9973 => x"81",
          9974 => x"81",
          9975 => x"7c",
          9976 => x"96",
          9977 => x"34",
          9978 => x"84",
          9979 => x"33",
          9980 => x"81",
          9981 => x"33",
          9982 => x"a4",
          9983 => x"e4",
          9984 => x"06",
          9985 => x"41",
          9986 => x"7f",
          9987 => x"78",
          9988 => x"38",
          9989 => x"81",
          9990 => x"58",
          9991 => x"38",
          9992 => x"83",
          9993 => x"0b",
          9994 => x"7a",
          9995 => x"81",
          9996 => x"b8",
          9997 => x"81",
          9998 => x"58",
          9999 => x"3f",
         10000 => x"08",
         10001 => x"38",
         10002 => x"59",
         10003 => x"0c",
         10004 => x"99",
         10005 => x"17",
         10006 => x"18",
         10007 => x"2b",
         10008 => x"83",
         10009 => x"d4",
         10010 => x"a5",
         10011 => x"26",
         10012 => x"b8",
         10013 => x"42",
         10014 => x"38",
         10015 => x"84",
         10016 => x"38",
         10017 => x"81",
         10018 => x"38",
         10019 => x"33",
         10020 => x"33",
         10021 => x"07",
         10022 => x"84",
         10023 => x"81",
         10024 => x"38",
         10025 => x"33",
         10026 => x"33",
         10027 => x"07",
         10028 => x"a4",
         10029 => x"17",
         10030 => x"82",
         10031 => x"90",
         10032 => x"2b",
         10033 => x"33",
         10034 => x"88",
         10035 => x"71",
         10036 => x"45",
         10037 => x"56",
         10038 => x"0c",
         10039 => x"33",
         10040 => x"80",
         10041 => x"ff",
         10042 => x"ff",
         10043 => x"59",
         10044 => x"81",
         10045 => x"38",
         10046 => x"06",
         10047 => x"80",
         10048 => x"5a",
         10049 => x"8a",
         10050 => x"59",
         10051 => x"87",
         10052 => x"18",
         10053 => x"61",
         10054 => x"80",
         10055 => x"80",
         10056 => x"71",
         10057 => x"56",
         10058 => x"18",
         10059 => x"8f",
         10060 => x"8d",
         10061 => x"98",
         10062 => x"17",
         10063 => x"18",
         10064 => x"2b",
         10065 => x"74",
         10066 => x"d8",
         10067 => x"33",
         10068 => x"71",
         10069 => x"88",
         10070 => x"14",
         10071 => x"07",
         10072 => x"33",
         10073 => x"44",
         10074 => x"42",
         10075 => x"17",
         10076 => x"18",
         10077 => x"2b",
         10078 => x"8d",
         10079 => x"2e",
         10080 => x"7d",
         10081 => x"2a",
         10082 => x"75",
         10083 => x"38",
         10084 => x"7a",
         10085 => x"ee",
         10086 => x"b8",
         10087 => x"84",
         10088 => x"80",
         10089 => x"38",
         10090 => x"08",
         10091 => x"ff",
         10092 => x"38",
         10093 => x"83",
         10094 => x"83",
         10095 => x"75",
         10096 => x"85",
         10097 => x"5d",
         10098 => x"9c",
         10099 => x"a4",
         10100 => x"1d",
         10101 => x"0c",
         10102 => x"1a",
         10103 => x"7c",
         10104 => x"87",
         10105 => x"22",
         10106 => x"7b",
         10107 => x"e0",
         10108 => x"ac",
         10109 => x"19",
         10110 => x"2e",
         10111 => x"10",
         10112 => x"2a",
         10113 => x"05",
         10114 => x"ff",
         10115 => x"59",
         10116 => x"a0",
         10117 => x"b8",
         10118 => x"94",
         10119 => x"0b",
         10120 => x"ff",
         10121 => x"18",
         10122 => x"2e",
         10123 => x"7c",
         10124 => x"d0",
         10125 => x"05",
         10126 => x"d0",
         10127 => x"86",
         10128 => x"d0",
         10129 => x"18",
         10130 => x"98",
         10131 => x"58",
         10132 => x"e4",
         10133 => x"0d",
         10134 => x"84",
         10135 => x"97",
         10136 => x"76",
         10137 => x"70",
         10138 => x"57",
         10139 => x"89",
         10140 => x"82",
         10141 => x"ff",
         10142 => x"5d",
         10143 => x"2e",
         10144 => x"80",
         10145 => x"e4",
         10146 => x"5c",
         10147 => x"5a",
         10148 => x"81",
         10149 => x"79",
         10150 => x"5b",
         10151 => x"12",
         10152 => x"77",
         10153 => x"38",
         10154 => x"81",
         10155 => x"55",
         10156 => x"58",
         10157 => x"89",
         10158 => x"70",
         10159 => x"58",
         10160 => x"70",
         10161 => x"55",
         10162 => x"09",
         10163 => x"38",
         10164 => x"38",
         10165 => x"70",
         10166 => x"07",
         10167 => x"07",
         10168 => x"7a",
         10169 => x"98",
         10170 => x"84",
         10171 => x"83",
         10172 => x"98",
         10173 => x"f9",
         10174 => x"80",
         10175 => x"38",
         10176 => x"81",
         10177 => x"58",
         10178 => x"38",
         10179 => x"c0",
         10180 => x"33",
         10181 => x"81",
         10182 => x"81",
         10183 => x"81",
         10184 => x"eb",
         10185 => x"70",
         10186 => x"07",
         10187 => x"77",
         10188 => x"75",
         10189 => x"83",
         10190 => x"3d",
         10191 => x"83",
         10192 => x"16",
         10193 => x"5b",
         10194 => x"a5",
         10195 => x"16",
         10196 => x"17",
         10197 => x"2b",
         10198 => x"07",
         10199 => x"33",
         10200 => x"88",
         10201 => x"1b",
         10202 => x"52",
         10203 => x"40",
         10204 => x"70",
         10205 => x"0c",
         10206 => x"17",
         10207 => x"80",
         10208 => x"38",
         10209 => x"1d",
         10210 => x"70",
         10211 => x"71",
         10212 => x"71",
         10213 => x"f0",
         10214 => x"1c",
         10215 => x"43",
         10216 => x"08",
         10217 => x"7a",
         10218 => x"fb",
         10219 => x"83",
         10220 => x"0b",
         10221 => x"7a",
         10222 => x"7a",
         10223 => x"38",
         10224 => x"53",
         10225 => x"81",
         10226 => x"ff",
         10227 => x"84",
         10228 => x"76",
         10229 => x"ff",
         10230 => x"74",
         10231 => x"84",
         10232 => x"38",
         10233 => x"7f",
         10234 => x"2b",
         10235 => x"83",
         10236 => x"d4",
         10237 => x"81",
         10238 => x"80",
         10239 => x"33",
         10240 => x"81",
         10241 => x"b7",
         10242 => x"eb",
         10243 => x"70",
         10244 => x"07",
         10245 => x"7f",
         10246 => x"81",
         10247 => x"38",
         10248 => x"81",
         10249 => x"80",
         10250 => x"d9",
         10251 => x"58",
         10252 => x"09",
         10253 => x"38",
         10254 => x"76",
         10255 => x"38",
         10256 => x"f8",
         10257 => x"1a",
         10258 => x"5a",
         10259 => x"fe",
         10260 => x"a8",
         10261 => x"80",
         10262 => x"e4",
         10263 => x"58",
         10264 => x"05",
         10265 => x"70",
         10266 => x"33",
         10267 => x"ff",
         10268 => x"56",
         10269 => x"2e",
         10270 => x"75",
         10271 => x"38",
         10272 => x"8a",
         10273 => x"98",
         10274 => x"7b",
         10275 => x"5d",
         10276 => x"81",
         10277 => x"71",
         10278 => x"1b",
         10279 => x"40",
         10280 => x"85",
         10281 => x"80",
         10282 => x"82",
         10283 => x"39",
         10284 => x"fa",
         10285 => x"84",
         10286 => x"97",
         10287 => x"75",
         10288 => x"2e",
         10289 => x"85",
         10290 => x"18",
         10291 => x"40",
         10292 => x"b7",
         10293 => x"84",
         10294 => x"97",
         10295 => x"83",
         10296 => x"18",
         10297 => x"5c",
         10298 => x"70",
         10299 => x"33",
         10300 => x"05",
         10301 => x"71",
         10302 => x"5b",
         10303 => x"77",
         10304 => x"d1",
         10305 => x"2e",
         10306 => x"0b",
         10307 => x"83",
         10308 => x"5a",
         10309 => x"81",
         10310 => x"7a",
         10311 => x"5c",
         10312 => x"31",
         10313 => x"58",
         10314 => x"80",
         10315 => x"38",
         10316 => x"e1",
         10317 => x"77",
         10318 => x"59",
         10319 => x"81",
         10320 => x"39",
         10321 => x"33",
         10322 => x"33",
         10323 => x"07",
         10324 => x"81",
         10325 => x"06",
         10326 => x"81",
         10327 => x"5a",
         10328 => x"78",
         10329 => x"83",
         10330 => x"7a",
         10331 => x"81",
         10332 => x"38",
         10333 => x"53",
         10334 => x"81",
         10335 => x"ff",
         10336 => x"84",
         10337 => x"80",
         10338 => x"ff",
         10339 => x"77",
         10340 => x"79",
         10341 => x"79",
         10342 => x"84",
         10343 => x"84",
         10344 => x"71",
         10345 => x"57",
         10346 => x"d4",
         10347 => x"81",
         10348 => x"38",
         10349 => x"11",
         10350 => x"33",
         10351 => x"71",
         10352 => x"81",
         10353 => x"72",
         10354 => x"75",
         10355 => x"5e",
         10356 => x"42",
         10357 => x"84",
         10358 => x"d2",
         10359 => x"06",
         10360 => x"84",
         10361 => x"11",
         10362 => x"33",
         10363 => x"71",
         10364 => x"81",
         10365 => x"72",
         10366 => x"75",
         10367 => x"47",
         10368 => x"5c",
         10369 => x"86",
         10370 => x"f2",
         10371 => x"06",
         10372 => x"84",
         10373 => x"11",
         10374 => x"33",
         10375 => x"71",
         10376 => x"81",
         10377 => x"72",
         10378 => x"75",
         10379 => x"94",
         10380 => x"84",
         10381 => x"11",
         10382 => x"33",
         10383 => x"71",
         10384 => x"81",
         10385 => x"72",
         10386 => x"75",
         10387 => x"62",
         10388 => x"59",
         10389 => x"5c",
         10390 => x"5b",
         10391 => x"77",
         10392 => x"bc",
         10393 => x"5d",
         10394 => x"bc",
         10395 => x"18",
         10396 => x"c4",
         10397 => x"0c",
         10398 => x"18",
         10399 => x"39",
         10400 => x"f8",
         10401 => x"7a",
         10402 => x"f2",
         10403 => x"54",
         10404 => x"53",
         10405 => x"53",
         10406 => x"52",
         10407 => x"b3",
         10408 => x"e4",
         10409 => x"09",
         10410 => x"a4",
         10411 => x"e4",
         10412 => x"34",
         10413 => x"a8",
         10414 => x"40",
         10415 => x"08",
         10416 => x"82",
         10417 => x"60",
         10418 => x"8d",
         10419 => x"e4",
         10420 => x"a0",
         10421 => x"74",
         10422 => x"91",
         10423 => x"81",
         10424 => x"e4",
         10425 => x"58",
         10426 => x"80",
         10427 => x"80",
         10428 => x"71",
         10429 => x"5f",
         10430 => x"7d",
         10431 => x"88",
         10432 => x"61",
         10433 => x"80",
         10434 => x"11",
         10435 => x"33",
         10436 => x"71",
         10437 => x"81",
         10438 => x"72",
         10439 => x"75",
         10440 => x"ac",
         10441 => x"7d",
         10442 => x"43",
         10443 => x"40",
         10444 => x"75",
         10445 => x"2e",
         10446 => x"82",
         10447 => x"39",
         10448 => x"f2",
         10449 => x"3d",
         10450 => x"83",
         10451 => x"39",
         10452 => x"f5",
         10453 => x"bf",
         10454 => x"b4",
         10455 => x"18",
         10456 => x"78",
         10457 => x"33",
         10458 => x"e7",
         10459 => x"39",
         10460 => x"02",
         10461 => x"33",
         10462 => x"93",
         10463 => x"5d",
         10464 => x"40",
         10465 => x"80",
         10466 => x"70",
         10467 => x"33",
         10468 => x"55",
         10469 => x"2e",
         10470 => x"73",
         10471 => x"ba",
         10472 => x"38",
         10473 => x"33",
         10474 => x"24",
         10475 => x"73",
         10476 => x"d0",
         10477 => x"08",
         10478 => x"80",
         10479 => x"80",
         10480 => x"54",
         10481 => x"86",
         10482 => x"34",
         10483 => x"75",
         10484 => x"7c",
         10485 => x"38",
         10486 => x"3d",
         10487 => x"05",
         10488 => x"3f",
         10489 => x"08",
         10490 => x"b8",
         10491 => x"3d",
         10492 => x"0b",
         10493 => x"0c",
         10494 => x"04",
         10495 => x"11",
         10496 => x"06",
         10497 => x"73",
         10498 => x"38",
         10499 => x"81",
         10500 => x"05",
         10501 => x"79",
         10502 => x"38",
         10503 => x"83",
         10504 => x"5f",
         10505 => x"7e",
         10506 => x"70",
         10507 => x"33",
         10508 => x"05",
         10509 => x"9f",
         10510 => x"55",
         10511 => x"89",
         10512 => x"70",
         10513 => x"56",
         10514 => x"16",
         10515 => x"26",
         10516 => x"16",
         10517 => x"06",
         10518 => x"30",
         10519 => x"58",
         10520 => x"2e",
         10521 => x"85",
         10522 => x"be",
         10523 => x"32",
         10524 => x"72",
         10525 => x"79",
         10526 => x"54",
         10527 => x"92",
         10528 => x"84",
         10529 => x"83",
         10530 => x"99",
         10531 => x"fe",
         10532 => x"83",
         10533 => x"7a",
         10534 => x"54",
         10535 => x"e6",
         10536 => x"02",
         10537 => x"fb",
         10538 => x"59",
         10539 => x"80",
         10540 => x"74",
         10541 => x"54",
         10542 => x"05",
         10543 => x"84",
         10544 => x"ed",
         10545 => x"b8",
         10546 => x"84",
         10547 => x"80",
         10548 => x"80",
         10549 => x"56",
         10550 => x"e4",
         10551 => x"0d",
         10552 => x"6d",
         10553 => x"70",
         10554 => x"9a",
         10555 => x"e4",
         10556 => x"b8",
         10557 => x"2e",
         10558 => x"77",
         10559 => x"7c",
         10560 => x"ca",
         10561 => x"2e",
         10562 => x"76",
         10563 => x"ea",
         10564 => x"07",
         10565 => x"bb",
         10566 => x"2a",
         10567 => x"7a",
         10568 => x"d1",
         10569 => x"11",
         10570 => x"33",
         10571 => x"07",
         10572 => x"42",
         10573 => x"56",
         10574 => x"84",
         10575 => x"0b",
         10576 => x"80",
         10577 => x"34",
         10578 => x"17",
         10579 => x"0b",
         10580 => x"66",
         10581 => x"8b",
         10582 => x"67",
         10583 => x"0b",
         10584 => x"80",
         10585 => x"34",
         10586 => x"7c",
         10587 => x"a9",
         10588 => x"80",
         10589 => x"34",
         10590 => x"1c",
         10591 => x"9e",
         10592 => x"0b",
         10593 => x"7e",
         10594 => x"83",
         10595 => x"80",
         10596 => x"38",
         10597 => x"08",
         10598 => x"53",
         10599 => x"81",
         10600 => x"38",
         10601 => x"7c",
         10602 => x"38",
         10603 => x"79",
         10604 => x"39",
         10605 => x"05",
         10606 => x"2b",
         10607 => x"80",
         10608 => x"38",
         10609 => x"06",
         10610 => x"fe",
         10611 => x"fe",
         10612 => x"80",
         10613 => x"70",
         10614 => x"06",
         10615 => x"82",
         10616 => x"81",
         10617 => x"5e",
         10618 => x"89",
         10619 => x"06",
         10620 => x"f6",
         10621 => x"2a",
         10622 => x"75",
         10623 => x"38",
         10624 => x"07",
         10625 => x"11",
         10626 => x"0c",
         10627 => x"0c",
         10628 => x"33",
         10629 => x"71",
         10630 => x"73",
         10631 => x"40",
         10632 => x"83",
         10633 => x"38",
         10634 => x"0c",
         10635 => x"11",
         10636 => x"33",
         10637 => x"71",
         10638 => x"81",
         10639 => x"72",
         10640 => x"75",
         10641 => x"70",
         10642 => x"0c",
         10643 => x"51",
         10644 => x"57",
         10645 => x"1a",
         10646 => x"23",
         10647 => x"34",
         10648 => x"1a",
         10649 => x"9c",
         10650 => x"85",
         10651 => x"55",
         10652 => x"84",
         10653 => x"80",
         10654 => x"38",
         10655 => x"0c",
         10656 => x"70",
         10657 => x"52",
         10658 => x"30",
         10659 => x"80",
         10660 => x"79",
         10661 => x"92",
         10662 => x"76",
         10663 => x"7d",
         10664 => x"86",
         10665 => x"78",
         10666 => x"db",
         10667 => x"e4",
         10668 => x"b8",
         10669 => x"26",
         10670 => x"57",
         10671 => x"08",
         10672 => x"cb",
         10673 => x"31",
         10674 => x"02",
         10675 => x"33",
         10676 => x"7d",
         10677 => x"82",
         10678 => x"55",
         10679 => x"fc",
         10680 => x"57",
         10681 => x"fb",
         10682 => x"57",
         10683 => x"fb",
         10684 => x"57",
         10685 => x"fb",
         10686 => x"51",
         10687 => x"84",
         10688 => x"78",
         10689 => x"57",
         10690 => x"38",
         10691 => x"7a",
         10692 => x"57",
         10693 => x"39",
         10694 => x"94",
         10695 => x"98",
         10696 => x"2b",
         10697 => x"5d",
         10698 => x"fc",
         10699 => x"7c",
         10700 => x"bd",
         10701 => x"79",
         10702 => x"cb",
         10703 => x"e4",
         10704 => x"b8",
         10705 => x"2e",
         10706 => x"84",
         10707 => x"81",
         10708 => x"38",
         10709 => x"08",
         10710 => x"99",
         10711 => x"74",
         10712 => x"ff",
         10713 => x"84",
         10714 => x"83",
         10715 => x"17",
         10716 => x"94",
         10717 => x"56",
         10718 => x"27",
         10719 => x"81",
         10720 => x"0c",
         10721 => x"81",
         10722 => x"84",
         10723 => x"55",
         10724 => x"ff",
         10725 => x"d9",
         10726 => x"94",
         10727 => x"0b",
         10728 => x"fb",
         10729 => x"16",
         10730 => x"33",
         10731 => x"71",
         10732 => x"7e",
         10733 => x"5b",
         10734 => x"17",
         10735 => x"8f",
         10736 => x"0b",
         10737 => x"80",
         10738 => x"17",
         10739 => x"a0",
         10740 => x"34",
         10741 => x"5e",
         10742 => x"17",
         10743 => x"9b",
         10744 => x"33",
         10745 => x"2e",
         10746 => x"fb",
         10747 => x"a9",
         10748 => x"7f",
         10749 => x"57",
         10750 => x"08",
         10751 => x"38",
         10752 => x"5a",
         10753 => x"09",
         10754 => x"38",
         10755 => x"53",
         10756 => x"81",
         10757 => x"ff",
         10758 => x"84",
         10759 => x"80",
         10760 => x"ff",
         10761 => x"76",
         10762 => x"7e",
         10763 => x"1d",
         10764 => x"57",
         10765 => x"fb",
         10766 => x"79",
         10767 => x"39",
         10768 => x"16",
         10769 => x"16",
         10770 => x"17",
         10771 => x"ff",
         10772 => x"84",
         10773 => x"7d",
         10774 => x"06",
         10775 => x"84",
         10776 => x"83",
         10777 => x"16",
         10778 => x"08",
         10779 => x"e4",
         10780 => x"74",
         10781 => x"27",
         10782 => x"82",
         10783 => x"74",
         10784 => x"81",
         10785 => x"38",
         10786 => x"16",
         10787 => x"08",
         10788 => x"52",
         10789 => x"51",
         10790 => x"3f",
         10791 => x"ec",
         10792 => x"1a",
         10793 => x"f8",
         10794 => x"98",
         10795 => x"f8",
         10796 => x"83",
         10797 => x"79",
         10798 => x"9a",
         10799 => x"19",
         10800 => x"fe",
         10801 => x"5a",
         10802 => x"f9",
         10803 => x"1a",
         10804 => x"29",
         10805 => x"05",
         10806 => x"80",
         10807 => x"38",
         10808 => x"15",
         10809 => x"76",
         10810 => x"39",
         10811 => x"0c",
         10812 => x"e4",
         10813 => x"80",
         10814 => x"da",
         10815 => x"e4",
         10816 => x"79",
         10817 => x"39",
         10818 => x"5b",
         10819 => x"f0",
         10820 => x"65",
         10821 => x"40",
         10822 => x"7e",
         10823 => x"79",
         10824 => x"38",
         10825 => x"75",
         10826 => x"38",
         10827 => x"74",
         10828 => x"38",
         10829 => x"84",
         10830 => x"59",
         10831 => x"84",
         10832 => x"55",
         10833 => x"55",
         10834 => x"38",
         10835 => x"55",
         10836 => x"38",
         10837 => x"81",
         10838 => x"56",
         10839 => x"81",
         10840 => x"1a",
         10841 => x"08",
         10842 => x"56",
         10843 => x"81",
         10844 => x"80",
         10845 => x"38",
         10846 => x"83",
         10847 => x"7a",
         10848 => x"8a",
         10849 => x"05",
         10850 => x"06",
         10851 => x"38",
         10852 => x"38",
         10853 => x"55",
         10854 => x"84",
         10855 => x"ff",
         10856 => x"38",
         10857 => x"0c",
         10858 => x"1a",
         10859 => x"9c",
         10860 => x"05",
         10861 => x"60",
         10862 => x"38",
         10863 => x"70",
         10864 => x"1b",
         10865 => x"56",
         10866 => x"83",
         10867 => x"15",
         10868 => x"59",
         10869 => x"2e",
         10870 => x"77",
         10871 => x"75",
         10872 => x"75",
         10873 => x"77",
         10874 => x"7c",
         10875 => x"33",
         10876 => x"e0",
         10877 => x"e4",
         10878 => x"38",
         10879 => x"33",
         10880 => x"80",
         10881 => x"b4",
         10882 => x"31",
         10883 => x"27",
         10884 => x"80",
         10885 => x"1e",
         10886 => x"58",
         10887 => x"81",
         10888 => x"77",
         10889 => x"59",
         10890 => x"55",
         10891 => x"77",
         10892 => x"7b",
         10893 => x"08",
         10894 => x"78",
         10895 => x"08",
         10896 => x"94",
         10897 => x"5c",
         10898 => x"38",
         10899 => x"84",
         10900 => x"92",
         10901 => x"74",
         10902 => x"0c",
         10903 => x"04",
         10904 => x"8e",
         10905 => x"08",
         10906 => x"ff",
         10907 => x"71",
         10908 => x"7b",
         10909 => x"38",
         10910 => x"56",
         10911 => x"77",
         10912 => x"80",
         10913 => x"33",
         10914 => x"5f",
         10915 => x"09",
         10916 => x"e4",
         10917 => x"76",
         10918 => x"52",
         10919 => x"51",
         10920 => x"3f",
         10921 => x"08",
         10922 => x"38",
         10923 => x"5b",
         10924 => x"0c",
         10925 => x"38",
         10926 => x"08",
         10927 => x"11",
         10928 => x"58",
         10929 => x"59",
         10930 => x"fe",
         10931 => x"70",
         10932 => x"33",
         10933 => x"05",
         10934 => x"16",
         10935 => x"2e",
         10936 => x"74",
         10937 => x"56",
         10938 => x"81",
         10939 => x"ff",
         10940 => x"da",
         10941 => x"39",
         10942 => x"19",
         10943 => x"19",
         10944 => x"1a",
         10945 => x"ff",
         10946 => x"81",
         10947 => x"e4",
         10948 => x"09",
         10949 => x"9c",
         10950 => x"e4",
         10951 => x"34",
         10952 => x"a8",
         10953 => x"84",
         10954 => x"5c",
         10955 => x"1a",
         10956 => x"e1",
         10957 => x"33",
         10958 => x"2e",
         10959 => x"fe",
         10960 => x"54",
         10961 => x"a0",
         10962 => x"53",
         10963 => x"19",
         10964 => x"9d",
         10965 => x"5b",
         10966 => x"76",
         10967 => x"94",
         10968 => x"fe",
         10969 => x"1a",
         10970 => x"51",
         10971 => x"3f",
         10972 => x"08",
         10973 => x"39",
         10974 => x"51",
         10975 => x"3f",
         10976 => x"08",
         10977 => x"74",
         10978 => x"74",
         10979 => x"57",
         10980 => x"81",
         10981 => x"34",
         10982 => x"b8",
         10983 => x"3d",
         10984 => x"0b",
         10985 => x"82",
         10986 => x"e4",
         10987 => x"0d",
         10988 => x"0d",
         10989 => x"66",
         10990 => x"5a",
         10991 => x"89",
         10992 => x"2e",
         10993 => x"08",
         10994 => x"2e",
         10995 => x"33",
         10996 => x"2e",
         10997 => x"16",
         10998 => x"22",
         10999 => x"78",
         11000 => x"38",
         11001 => x"41",
         11002 => x"82",
         11003 => x"1a",
         11004 => x"82",
         11005 => x"1a",
         11006 => x"2a",
         11007 => x"58",
         11008 => x"80",
         11009 => x"38",
         11010 => x"7b",
         11011 => x"7b",
         11012 => x"38",
         11013 => x"7a",
         11014 => x"81",
         11015 => x"ff",
         11016 => x"82",
         11017 => x"8a",
         11018 => x"05",
         11019 => x"06",
         11020 => x"aa",
         11021 => x"9e",
         11022 => x"08",
         11023 => x"2e",
         11024 => x"74",
         11025 => x"a1",
         11026 => x"2e",
         11027 => x"74",
         11028 => x"88",
         11029 => x"38",
         11030 => x"0c",
         11031 => x"16",
         11032 => x"08",
         11033 => x"38",
         11034 => x"fe",
         11035 => x"08",
         11036 => x"58",
         11037 => x"85",
         11038 => x"16",
         11039 => x"29",
         11040 => x"05",
         11041 => x"80",
         11042 => x"38",
         11043 => x"89",
         11044 => x"77",
         11045 => x"98",
         11046 => x"5f",
         11047 => x"85",
         11048 => x"31",
         11049 => x"7b",
         11050 => x"81",
         11051 => x"ff",
         11052 => x"84",
         11053 => x"85",
         11054 => x"b4",
         11055 => x"31",
         11056 => x"78",
         11057 => x"84",
         11058 => x"18",
         11059 => x"1f",
         11060 => x"74",
         11061 => x"56",
         11062 => x"81",
         11063 => x"ff",
         11064 => x"ef",
         11065 => x"75",
         11066 => x"77",
         11067 => x"7a",
         11068 => x"08",
         11069 => x"79",
         11070 => x"08",
         11071 => x"94",
         11072 => x"1e",
         11073 => x"57",
         11074 => x"75",
         11075 => x"74",
         11076 => x"1b",
         11077 => x"85",
         11078 => x"33",
         11079 => x"c0",
         11080 => x"90",
         11081 => x"56",
         11082 => x"e4",
         11083 => x"0d",
         11084 => x"b8",
         11085 => x"3d",
         11086 => x"16",
         11087 => x"82",
         11088 => x"56",
         11089 => x"60",
         11090 => x"59",
         11091 => x"ff",
         11092 => x"71",
         11093 => x"7a",
         11094 => x"38",
         11095 => x"57",
         11096 => x"78",
         11097 => x"80",
         11098 => x"33",
         11099 => x"5f",
         11100 => x"09",
         11101 => x"d5",
         11102 => x"77",
         11103 => x"52",
         11104 => x"51",
         11105 => x"3f",
         11106 => x"08",
         11107 => x"38",
         11108 => x"5c",
         11109 => x"0c",
         11110 => x"38",
         11111 => x"08",
         11112 => x"11",
         11113 => x"05",
         11114 => x"58",
         11115 => x"95",
         11116 => x"81",
         11117 => x"75",
         11118 => x"57",
         11119 => x"56",
         11120 => x"60",
         11121 => x"83",
         11122 => x"a3",
         11123 => x"b4",
         11124 => x"b8",
         11125 => x"81",
         11126 => x"40",
         11127 => x"3f",
         11128 => x"b8",
         11129 => x"2e",
         11130 => x"ff",
         11131 => x"b8",
         11132 => x"17",
         11133 => x"08",
         11134 => x"31",
         11135 => x"08",
         11136 => x"a0",
         11137 => x"fe",
         11138 => x"16",
         11139 => x"82",
         11140 => x"06",
         11141 => x"81",
         11142 => x"08",
         11143 => x"05",
         11144 => x"81",
         11145 => x"ff",
         11146 => x"7e",
         11147 => x"39",
         11148 => x"57",
         11149 => x"77",
         11150 => x"83",
         11151 => x"7f",
         11152 => x"60",
         11153 => x"0c",
         11154 => x"58",
         11155 => x"9c",
         11156 => x"fd",
         11157 => x"1a",
         11158 => x"51",
         11159 => x"3f",
         11160 => x"08",
         11161 => x"e4",
         11162 => x"38",
         11163 => x"58",
         11164 => x"76",
         11165 => x"ff",
         11166 => x"84",
         11167 => x"55",
         11168 => x"08",
         11169 => x"e4",
         11170 => x"b4",
         11171 => x"b8",
         11172 => x"81",
         11173 => x"57",
         11174 => x"3f",
         11175 => x"08",
         11176 => x"84",
         11177 => x"83",
         11178 => x"16",
         11179 => x"08",
         11180 => x"a0",
         11181 => x"fd",
         11182 => x"16",
         11183 => x"82",
         11184 => x"06",
         11185 => x"81",
         11186 => x"08",
         11187 => x"05",
         11188 => x"81",
         11189 => x"ff",
         11190 => x"60",
         11191 => x"39",
         11192 => x"51",
         11193 => x"3f",
         11194 => x"08",
         11195 => x"74",
         11196 => x"74",
         11197 => x"57",
         11198 => x"81",
         11199 => x"08",
         11200 => x"70",
         11201 => x"33",
         11202 => x"96",
         11203 => x"b8",
         11204 => x"c6",
         11205 => x"e4",
         11206 => x"34",
         11207 => x"a8",
         11208 => x"55",
         11209 => x"08",
         11210 => x"38",
         11211 => x"58",
         11212 => x"09",
         11213 => x"8b",
         11214 => x"b4",
         11215 => x"17",
         11216 => x"76",
         11217 => x"33",
         11218 => x"87",
         11219 => x"b4",
         11220 => x"1b",
         11221 => x"fd",
         11222 => x"0b",
         11223 => x"81",
         11224 => x"e4",
         11225 => x"0d",
         11226 => x"91",
         11227 => x"0b",
         11228 => x"0c",
         11229 => x"04",
         11230 => x"7d",
         11231 => x"77",
         11232 => x"38",
         11233 => x"75",
         11234 => x"38",
         11235 => x"74",
         11236 => x"38",
         11237 => x"84",
         11238 => x"59",
         11239 => x"83",
         11240 => x"55",
         11241 => x"56",
         11242 => x"38",
         11243 => x"70",
         11244 => x"06",
         11245 => x"80",
         11246 => x"38",
         11247 => x"08",
         11248 => x"17",
         11249 => x"ac",
         11250 => x"33",
         11251 => x"bc",
         11252 => x"78",
         11253 => x"52",
         11254 => x"51",
         11255 => x"3f",
         11256 => x"08",
         11257 => x"38",
         11258 => x"56",
         11259 => x"0c",
         11260 => x"38",
         11261 => x"8b",
         11262 => x"07",
         11263 => x"8b",
         11264 => x"08",
         11265 => x"70",
         11266 => x"06",
         11267 => x"7a",
         11268 => x"7a",
         11269 => x"79",
         11270 => x"9c",
         11271 => x"96",
         11272 => x"5b",
         11273 => x"81",
         11274 => x"18",
         11275 => x"7b",
         11276 => x"2a",
         11277 => x"18",
         11278 => x"2a",
         11279 => x"18",
         11280 => x"2a",
         11281 => x"18",
         11282 => x"34",
         11283 => x"18",
         11284 => x"98",
         11285 => x"cc",
         11286 => x"34",
         11287 => x"18",
         11288 => x"93",
         11289 => x"5b",
         11290 => x"1c",
         11291 => x"ff",
         11292 => x"84",
         11293 => x"90",
         11294 => x"bf",
         11295 => x"79",
         11296 => x"75",
         11297 => x"0c",
         11298 => x"04",
         11299 => x"17",
         11300 => x"17",
         11301 => x"18",
         11302 => x"ff",
         11303 => x"81",
         11304 => x"e4",
         11305 => x"38",
         11306 => x"08",
         11307 => x"b4",
         11308 => x"18",
         11309 => x"b8",
         11310 => x"55",
         11311 => x"08",
         11312 => x"38",
         11313 => x"55",
         11314 => x"09",
         11315 => x"81",
         11316 => x"b4",
         11317 => x"18",
         11318 => x"7a",
         11319 => x"33",
         11320 => x"ef",
         11321 => x"fd",
         11322 => x"90",
         11323 => x"94",
         11324 => x"88",
         11325 => x"95",
         11326 => x"18",
         11327 => x"7b",
         11328 => x"2a",
         11329 => x"18",
         11330 => x"2a",
         11331 => x"18",
         11332 => x"2a",
         11333 => x"18",
         11334 => x"34",
         11335 => x"18",
         11336 => x"98",
         11337 => x"cc",
         11338 => x"34",
         11339 => x"18",
         11340 => x"93",
         11341 => x"5b",
         11342 => x"1c",
         11343 => x"ff",
         11344 => x"84",
         11345 => x"90",
         11346 => x"bf",
         11347 => x"79",
         11348 => x"fe",
         11349 => x"16",
         11350 => x"90",
         11351 => x"b8",
         11352 => x"06",
         11353 => x"ba",
         11354 => x"08",
         11355 => x"b4",
         11356 => x"0d",
         11357 => x"55",
         11358 => x"84",
         11359 => x"54",
         11360 => x"08",
         11361 => x"56",
         11362 => x"9e",
         11363 => x"53",
         11364 => x"96",
         11365 => x"52",
         11366 => x"8e",
         11367 => x"22",
         11368 => x"58",
         11369 => x"2e",
         11370 => x"52",
         11371 => x"54",
         11372 => x"75",
         11373 => x"84",
         11374 => x"89",
         11375 => x"81",
         11376 => x"ff",
         11377 => x"84",
         11378 => x"81",
         11379 => x"da",
         11380 => x"08",
         11381 => x"39",
         11382 => x"ff",
         11383 => x"57",
         11384 => x"2e",
         11385 => x"70",
         11386 => x"33",
         11387 => x"52",
         11388 => x"2e",
         11389 => x"ee",
         11390 => x"2e",
         11391 => x"d0",
         11392 => x"80",
         11393 => x"38",
         11394 => x"c0",
         11395 => x"84",
         11396 => x"8c",
         11397 => x"8b",
         11398 => x"e4",
         11399 => x"0d",
         11400 => x"d0",
         11401 => x"ff",
         11402 => x"53",
         11403 => x"91",
         11404 => x"73",
         11405 => x"d0",
         11406 => x"73",
         11407 => x"f5",
         11408 => x"83",
         11409 => x"58",
         11410 => x"56",
         11411 => x"81",
         11412 => x"75",
         11413 => x"57",
         11414 => x"12",
         11415 => x"70",
         11416 => x"38",
         11417 => x"81",
         11418 => x"54",
         11419 => x"51",
         11420 => x"89",
         11421 => x"70",
         11422 => x"54",
         11423 => x"70",
         11424 => x"51",
         11425 => x"09",
         11426 => x"38",
         11427 => x"38",
         11428 => x"70",
         11429 => x"07",
         11430 => x"07",
         11431 => x"76",
         11432 => x"38",
         11433 => x"1b",
         11434 => x"78",
         11435 => x"38",
         11436 => x"cf",
         11437 => x"24",
         11438 => x"76",
         11439 => x"c3",
         11440 => x"0d",
         11441 => x"3d",
         11442 => x"99",
         11443 => x"94",
         11444 => x"e4",
         11445 => x"b8",
         11446 => x"2e",
         11447 => x"84",
         11448 => x"98",
         11449 => x"7a",
         11450 => x"98",
         11451 => x"51",
         11452 => x"84",
         11453 => x"55",
         11454 => x"08",
         11455 => x"02",
         11456 => x"33",
         11457 => x"58",
         11458 => x"24",
         11459 => x"02",
         11460 => x"70",
         11461 => x"06",
         11462 => x"80",
         11463 => x"7a",
         11464 => x"33",
         11465 => x"71",
         11466 => x"73",
         11467 => x"5b",
         11468 => x"83",
         11469 => x"76",
         11470 => x"74",
         11471 => x"0c",
         11472 => x"04",
         11473 => x"08",
         11474 => x"81",
         11475 => x"38",
         11476 => x"b8",
         11477 => x"3d",
         11478 => x"16",
         11479 => x"33",
         11480 => x"71",
         11481 => x"79",
         11482 => x"0c",
         11483 => x"39",
         11484 => x"12",
         11485 => x"84",
         11486 => x"98",
         11487 => x"ff",
         11488 => x"80",
         11489 => x"80",
         11490 => x"5d",
         11491 => x"34",
         11492 => x"e4",
         11493 => x"05",
         11494 => x"3d",
         11495 => x"3f",
         11496 => x"08",
         11497 => x"e4",
         11498 => x"38",
         11499 => x"3d",
         11500 => x"98",
         11501 => x"dd",
         11502 => x"80",
         11503 => x"5b",
         11504 => x"2e",
         11505 => x"80",
         11506 => x"3d",
         11507 => x"52",
         11508 => x"a4",
         11509 => x"b8",
         11510 => x"84",
         11511 => x"83",
         11512 => x"80",
         11513 => x"58",
         11514 => x"08",
         11515 => x"38",
         11516 => x"08",
         11517 => x"5f",
         11518 => x"c7",
         11519 => x"76",
         11520 => x"52",
         11521 => x"51",
         11522 => x"3f",
         11523 => x"08",
         11524 => x"38",
         11525 => x"59",
         11526 => x"0c",
         11527 => x"38",
         11528 => x"08",
         11529 => x"9a",
         11530 => x"88",
         11531 => x"70",
         11532 => x"59",
         11533 => x"83",
         11534 => x"38",
         11535 => x"3d",
         11536 => x"7a",
         11537 => x"b7",
         11538 => x"e4",
         11539 => x"b8",
         11540 => x"9f",
         11541 => x"7a",
         11542 => x"f5",
         11543 => x"e4",
         11544 => x"b8",
         11545 => x"38",
         11546 => x"08",
         11547 => x"9a",
         11548 => x"88",
         11549 => x"70",
         11550 => x"59",
         11551 => x"83",
         11552 => x"38",
         11553 => x"a4",
         11554 => x"e4",
         11555 => x"51",
         11556 => x"3f",
         11557 => x"08",
         11558 => x"e4",
         11559 => x"ff",
         11560 => x"84",
         11561 => x"38",
         11562 => x"38",
         11563 => x"fd",
         11564 => x"7a",
         11565 => x"89",
         11566 => x"82",
         11567 => x"57",
         11568 => x"90",
         11569 => x"56",
         11570 => x"17",
         11571 => x"57",
         11572 => x"38",
         11573 => x"75",
         11574 => x"95",
         11575 => x"2e",
         11576 => x"17",
         11577 => x"ff",
         11578 => x"3d",
         11579 => x"19",
         11580 => x"59",
         11581 => x"33",
         11582 => x"eb",
         11583 => x"80",
         11584 => x"11",
         11585 => x"7e",
         11586 => x"3d",
         11587 => x"fd",
         11588 => x"60",
         11589 => x"38",
         11590 => x"d0",
         11591 => x"10",
         11592 => x"d4",
         11593 => x"70",
         11594 => x"59",
         11595 => x"7a",
         11596 => x"81",
         11597 => x"70",
         11598 => x"5a",
         11599 => x"82",
         11600 => x"78",
         11601 => x"80",
         11602 => x"27",
         11603 => x"16",
         11604 => x"7c",
         11605 => x"5e",
         11606 => x"57",
         11607 => x"ee",
         11608 => x"70",
         11609 => x"34",
         11610 => x"09",
         11611 => x"df",
         11612 => x"80",
         11613 => x"84",
         11614 => x"80",
         11615 => x"04",
         11616 => x"94",
         11617 => x"98",
         11618 => x"2b",
         11619 => x"59",
         11620 => x"f0",
         11621 => x"33",
         11622 => x"71",
         11623 => x"90",
         11624 => x"07",
         11625 => x"0c",
         11626 => x"52",
         11627 => x"a0",
         11628 => x"b8",
         11629 => x"84",
         11630 => x"80",
         11631 => x"38",
         11632 => x"81",
         11633 => x"08",
         11634 => x"70",
         11635 => x"33",
         11636 => x"88",
         11637 => x"59",
         11638 => x"08",
         11639 => x"84",
         11640 => x"83",
         11641 => x"16",
         11642 => x"08",
         11643 => x"e4",
         11644 => x"74",
         11645 => x"27",
         11646 => x"82",
         11647 => x"74",
         11648 => x"81",
         11649 => x"38",
         11650 => x"16",
         11651 => x"08",
         11652 => x"52",
         11653 => x"51",
         11654 => x"3f",
         11655 => x"dd",
         11656 => x"80",
         11657 => x"11",
         11658 => x"7b",
         11659 => x"84",
         11660 => x"70",
         11661 => x"e4",
         11662 => x"08",
         11663 => x"59",
         11664 => x"7e",
         11665 => x"81",
         11666 => x"38",
         11667 => x"80",
         11668 => x"18",
         11669 => x"5a",
         11670 => x"70",
         11671 => x"34",
         11672 => x"fe",
         11673 => x"e5",
         11674 => x"81",
         11675 => x"79",
         11676 => x"81",
         11677 => x"7f",
         11678 => x"38",
         11679 => x"82",
         11680 => x"34",
         11681 => x"e4",
         11682 => x"3d",
         11683 => x"3d",
         11684 => x"58",
         11685 => x"74",
         11686 => x"38",
         11687 => x"73",
         11688 => x"38",
         11689 => x"72",
         11690 => x"38",
         11691 => x"84",
         11692 => x"59",
         11693 => x"83",
         11694 => x"53",
         11695 => x"53",
         11696 => x"38",
         11697 => x"53",
         11698 => x"38",
         11699 => x"56",
         11700 => x"81",
         11701 => x"15",
         11702 => x"58",
         11703 => x"81",
         11704 => x"8a",
         11705 => x"89",
         11706 => x"56",
         11707 => x"81",
         11708 => x"52",
         11709 => x"fd",
         11710 => x"84",
         11711 => x"ff",
         11712 => x"70",
         11713 => x"fd",
         11714 => x"84",
         11715 => x"73",
         11716 => x"38",
         11717 => x"06",
         11718 => x"0c",
         11719 => x"98",
         11720 => x"58",
         11721 => x"2e",
         11722 => x"75",
         11723 => x"d9",
         11724 => x"31",
         11725 => x"17",
         11726 => x"90",
         11727 => x"81",
         11728 => x"51",
         11729 => x"80",
         11730 => x"38",
         11731 => x"51",
         11732 => x"3f",
         11733 => x"08",
         11734 => x"e4",
         11735 => x"81",
         11736 => x"ff",
         11737 => x"81",
         11738 => x"b4",
         11739 => x"73",
         11740 => x"27",
         11741 => x"73",
         11742 => x"ff",
         11743 => x"0b",
         11744 => x"81",
         11745 => x"b8",
         11746 => x"3d",
         11747 => x"15",
         11748 => x"2a",
         11749 => x"58",
         11750 => x"38",
         11751 => x"08",
         11752 => x"58",
         11753 => x"09",
         11754 => x"b6",
         11755 => x"16",
         11756 => x"08",
         11757 => x"27",
         11758 => x"8c",
         11759 => x"15",
         11760 => x"07",
         11761 => x"16",
         11762 => x"ff",
         11763 => x"80",
         11764 => x"9c",
         11765 => x"2e",
         11766 => x"9c",
         11767 => x"0b",
         11768 => x"0c",
         11769 => x"04",
         11770 => x"16",
         11771 => x"08",
         11772 => x"2e",
         11773 => x"73",
         11774 => x"73",
         11775 => x"c2",
         11776 => x"39",
         11777 => x"08",
         11778 => x"08",
         11779 => x"0c",
         11780 => x"06",
         11781 => x"2e",
         11782 => x"fe",
         11783 => x"08",
         11784 => x"55",
         11785 => x"27",
         11786 => x"8a",
         11787 => x"71",
         11788 => x"08",
         11789 => x"2a",
         11790 => x"53",
         11791 => x"80",
         11792 => x"15",
         11793 => x"e9",
         11794 => x"74",
         11795 => x"b7",
         11796 => x"e4",
         11797 => x"8a",
         11798 => x"33",
         11799 => x"a2",
         11800 => x"e4",
         11801 => x"53",
         11802 => x"38",
         11803 => x"54",
         11804 => x"39",
         11805 => x"51",
         11806 => x"3f",
         11807 => x"08",
         11808 => x"e4",
         11809 => x"98",
         11810 => x"e4",
         11811 => x"fd",
         11812 => x"b8",
         11813 => x"16",
         11814 => x"16",
         11815 => x"39",
         11816 => x"16",
         11817 => x"84",
         11818 => x"8b",
         11819 => x"f6",
         11820 => x"56",
         11821 => x"80",
         11822 => x"80",
         11823 => x"fc",
         11824 => x"3d",
         11825 => x"c5",
         11826 => x"b8",
         11827 => x"84",
         11828 => x"80",
         11829 => x"80",
         11830 => x"54",
         11831 => x"e4",
         11832 => x"0d",
         11833 => x"0c",
         11834 => x"51",
         11835 => x"3f",
         11836 => x"08",
         11837 => x"e4",
         11838 => x"38",
         11839 => x"70",
         11840 => x"59",
         11841 => x"af",
         11842 => x"33",
         11843 => x"81",
         11844 => x"79",
         11845 => x"c5",
         11846 => x"08",
         11847 => x"9a",
         11848 => x"88",
         11849 => x"70",
         11850 => x"5a",
         11851 => x"83",
         11852 => x"77",
         11853 => x"7a",
         11854 => x"22",
         11855 => x"74",
         11856 => x"ff",
         11857 => x"84",
         11858 => x"55",
         11859 => x"8d",
         11860 => x"2e",
         11861 => x"80",
         11862 => x"fe",
         11863 => x"80",
         11864 => x"f6",
         11865 => x"33",
         11866 => x"71",
         11867 => x"90",
         11868 => x"07",
         11869 => x"5a",
         11870 => x"39",
         11871 => x"78",
         11872 => x"74",
         11873 => x"38",
         11874 => x"72",
         11875 => x"38",
         11876 => x"71",
         11877 => x"38",
         11878 => x"84",
         11879 => x"52",
         11880 => x"94",
         11881 => x"71",
         11882 => x"38",
         11883 => x"73",
         11884 => x"0c",
         11885 => x"04",
         11886 => x"51",
         11887 => x"3f",
         11888 => x"08",
         11889 => x"71",
         11890 => x"75",
         11891 => x"d7",
         11892 => x"0d",
         11893 => x"55",
         11894 => x"80",
         11895 => x"74",
         11896 => x"80",
         11897 => x"73",
         11898 => x"80",
         11899 => x"86",
         11900 => x"16",
         11901 => x"72",
         11902 => x"97",
         11903 => x"72",
         11904 => x"75",
         11905 => x"76",
         11906 => x"f3",
         11907 => x"74",
         11908 => x"bd",
         11909 => x"e4",
         11910 => x"b8",
         11911 => x"2e",
         11912 => x"b8",
         11913 => x"38",
         11914 => x"51",
         11915 => x"3f",
         11916 => x"51",
         11917 => x"3f",
         11918 => x"08",
         11919 => x"30",
         11920 => x"9f",
         11921 => x"e4",
         11922 => x"57",
         11923 => x"b8",
         11924 => x"3d",
         11925 => x"77",
         11926 => x"53",
         11927 => x"3f",
         11928 => x"51",
         11929 => x"3f",
         11930 => x"08",
         11931 => x"30",
         11932 => x"9f",
         11933 => x"e4",
         11934 => x"57",
         11935 => x"75",
         11936 => x"ff",
         11937 => x"84",
         11938 => x"84",
         11939 => x"8a",
         11940 => x"81",
         11941 => x"fe",
         11942 => x"84",
         11943 => x"81",
         11944 => x"fe",
         11945 => x"75",
         11946 => x"fe",
         11947 => x"3d",
         11948 => x"80",
         11949 => x"70",
         11950 => x"52",
         11951 => x"3f",
         11952 => x"08",
         11953 => x"e4",
         11954 => x"8a",
         11955 => x"b8",
         11956 => x"3d",
         11957 => x"52",
         11958 => x"b5",
         11959 => x"b8",
         11960 => x"84",
         11961 => x"e5",
         11962 => x"cb",
         11963 => x"98",
         11964 => x"80",
         11965 => x"38",
         11966 => x"d1",
         11967 => x"75",
         11968 => x"bd",
         11969 => x"b8",
         11970 => x"3d",
         11971 => x"0b",
         11972 => x"0c",
         11973 => x"04",
         11974 => x"66",
         11975 => x"80",
         11976 => x"ec",
         11977 => x"3d",
         11978 => x"3f",
         11979 => x"08",
         11980 => x"e4",
         11981 => x"7f",
         11982 => x"08",
         11983 => x"fe",
         11984 => x"08",
         11985 => x"57",
         11986 => x"8d",
         11987 => x"0c",
         11988 => x"e4",
         11989 => x"0d",
         11990 => x"e4",
         11991 => x"5a",
         11992 => x"2e",
         11993 => x"77",
         11994 => x"84",
         11995 => x"5a",
         11996 => x"80",
         11997 => x"81",
         11998 => x"5d",
         11999 => x"08",
         12000 => x"ef",
         12001 => x"33",
         12002 => x"7c",
         12003 => x"81",
         12004 => x"b8",
         12005 => x"17",
         12006 => x"fc",
         12007 => x"b8",
         12008 => x"2e",
         12009 => x"5a",
         12010 => x"b4",
         12011 => x"7e",
         12012 => x"80",
         12013 => x"33",
         12014 => x"2e",
         12015 => x"77",
         12016 => x"83",
         12017 => x"12",
         12018 => x"2b",
         12019 => x"07",
         12020 => x"70",
         12021 => x"2b",
         12022 => x"80",
         12023 => x"80",
         12024 => x"30",
         12025 => x"63",
         12026 => x"05",
         12027 => x"62",
         12028 => x"41",
         12029 => x"52",
         12030 => x"5e",
         12031 => x"f2",
         12032 => x"0c",
         12033 => x"0c",
         12034 => x"81",
         12035 => x"84",
         12036 => x"84",
         12037 => x"95",
         12038 => x"81",
         12039 => x"08",
         12040 => x"70",
         12041 => x"33",
         12042 => x"fc",
         12043 => x"5e",
         12044 => x"08",
         12045 => x"84",
         12046 => x"83",
         12047 => x"17",
         12048 => x"08",
         12049 => x"e4",
         12050 => x"74",
         12051 => x"27",
         12052 => x"82",
         12053 => x"74",
         12054 => x"81",
         12055 => x"38",
         12056 => x"17",
         12057 => x"08",
         12058 => x"52",
         12059 => x"51",
         12060 => x"3f",
         12061 => x"97",
         12062 => x"42",
         12063 => x"56",
         12064 => x"51",
         12065 => x"3f",
         12066 => x"08",
         12067 => x"e8",
         12068 => x"e4",
         12069 => x"80",
         12070 => x"b8",
         12071 => x"70",
         12072 => x"08",
         12073 => x"7c",
         12074 => x"62",
         12075 => x"5c",
         12076 => x"76",
         12077 => x"7a",
         12078 => x"94",
         12079 => x"17",
         12080 => x"58",
         12081 => x"34",
         12082 => x"77",
         12083 => x"81",
         12084 => x"33",
         12085 => x"07",
         12086 => x"80",
         12087 => x"1d",
         12088 => x"ff",
         12089 => x"5f",
         12090 => x"55",
         12091 => x"38",
         12092 => x"77",
         12093 => x"39",
         12094 => x"5a",
         12095 => x"7a",
         12096 => x"84",
         12097 => x"07",
         12098 => x"18",
         12099 => x"39",
         12100 => x"5a",
         12101 => x"3d",
         12102 => x"89",
         12103 => x"2e",
         12104 => x"08",
         12105 => x"2e",
         12106 => x"33",
         12107 => x"2e",
         12108 => x"15",
         12109 => x"22",
         12110 => x"78",
         12111 => x"38",
         12112 => x"5a",
         12113 => x"38",
         12114 => x"56",
         12115 => x"38",
         12116 => x"70",
         12117 => x"06",
         12118 => x"55",
         12119 => x"80",
         12120 => x"17",
         12121 => x"8c",
         12122 => x"b7",
         12123 => x"d5",
         12124 => x"08",
         12125 => x"54",
         12126 => x"88",
         12127 => x"08",
         12128 => x"38",
         12129 => x"0b",
         12130 => x"94",
         12131 => x"18",
         12132 => x"c0",
         12133 => x"90",
         12134 => x"80",
         12135 => x"75",
         12136 => x"75",
         12137 => x"b8",
         12138 => x"3d",
         12139 => x"54",
         12140 => x"80",
         12141 => x"52",
         12142 => x"fe",
         12143 => x"b8",
         12144 => x"84",
         12145 => x"80",
         12146 => x"38",
         12147 => x"08",
         12148 => x"d8",
         12149 => x"e4",
         12150 => x"82",
         12151 => x"53",
         12152 => x"51",
         12153 => x"3f",
         12154 => x"08",
         12155 => x"9c",
         12156 => x"11",
         12157 => x"57",
         12158 => x"74",
         12159 => x"38",
         12160 => x"17",
         12161 => x"33",
         12162 => x"73",
         12163 => x"78",
         12164 => x"26",
         12165 => x"9c",
         12166 => x"33",
         12167 => x"e2",
         12168 => x"e4",
         12169 => x"54",
         12170 => x"38",
         12171 => x"55",
         12172 => x"39",
         12173 => x"18",
         12174 => x"73",
         12175 => x"88",
         12176 => x"c7",
         12177 => x"08",
         12178 => x"fe",
         12179 => x"84",
         12180 => x"ff",
         12181 => x"38",
         12182 => x"08",
         12183 => x"be",
         12184 => x"ae",
         12185 => x"84",
         12186 => x"9c",
         12187 => x"81",
         12188 => x"b8",
         12189 => x"18",
         12190 => x"58",
         12191 => x"0b",
         12192 => x"08",
         12193 => x"38",
         12194 => x"08",
         12195 => x"27",
         12196 => x"74",
         12197 => x"38",
         12198 => x"52",
         12199 => x"83",
         12200 => x"b8",
         12201 => x"84",
         12202 => x"80",
         12203 => x"52",
         12204 => x"fc",
         12205 => x"b8",
         12206 => x"84",
         12207 => x"80",
         12208 => x"38",
         12209 => x"08",
         12210 => x"dc",
         12211 => x"e4",
         12212 => x"80",
         12213 => x"53",
         12214 => x"51",
         12215 => x"3f",
         12216 => x"08",
         12217 => x"9c",
         12218 => x"11",
         12219 => x"57",
         12220 => x"74",
         12221 => x"81",
         12222 => x"0c",
         12223 => x"81",
         12224 => x"84",
         12225 => x"54",
         12226 => x"ff",
         12227 => x"55",
         12228 => x"17",
         12229 => x"f3",
         12230 => x"fe",
         12231 => x"0b",
         12232 => x"59",
         12233 => x"39",
         12234 => x"39",
         12235 => x"18",
         12236 => x"fe",
         12237 => x"b8",
         12238 => x"18",
         12239 => x"fd",
         12240 => x"0b",
         12241 => x"59",
         12242 => x"39",
         12243 => x"08",
         12244 => x"81",
         12245 => x"39",
         12246 => x"82",
         12247 => x"ff",
         12248 => x"a8",
         12249 => x"b7",
         12250 => x"b8",
         12251 => x"84",
         12252 => x"80",
         12253 => x"75",
         12254 => x"0c",
         12255 => x"04",
         12256 => x"3d",
         12257 => x"3d",
         12258 => x"ff",
         12259 => x"84",
         12260 => x"56",
         12261 => x"08",
         12262 => x"81",
         12263 => x"70",
         12264 => x"06",
         12265 => x"56",
         12266 => x"76",
         12267 => x"80",
         12268 => x"38",
         12269 => x"05",
         12270 => x"06",
         12271 => x"56",
         12272 => x"38",
         12273 => x"08",
         12274 => x"9a",
         12275 => x"88",
         12276 => x"33",
         12277 => x"57",
         12278 => x"2e",
         12279 => x"76",
         12280 => x"06",
         12281 => x"2e",
         12282 => x"87",
         12283 => x"08",
         12284 => x"83",
         12285 => x"7a",
         12286 => x"e4",
         12287 => x"3d",
         12288 => x"ff",
         12289 => x"84",
         12290 => x"56",
         12291 => x"08",
         12292 => x"84",
         12293 => x"52",
         12294 => x"91",
         12295 => x"b8",
         12296 => x"84",
         12297 => x"a0",
         12298 => x"84",
         12299 => x"a7",
         12300 => x"95",
         12301 => x"17",
         12302 => x"2b",
         12303 => x"07",
         12304 => x"5d",
         12305 => x"39",
         12306 => x"08",
         12307 => x"38",
         12308 => x"08",
         12309 => x"78",
         12310 => x"3d",
         12311 => x"57",
         12312 => x"80",
         12313 => x"52",
         12314 => x"8b",
         12315 => x"b8",
         12316 => x"84",
         12317 => x"80",
         12318 => x"75",
         12319 => x"07",
         12320 => x"5a",
         12321 => x"9a",
         12322 => x"2e",
         12323 => x"79",
         12324 => x"81",
         12325 => x"38",
         12326 => x"7b",
         12327 => x"38",
         12328 => x"fd",
         12329 => x"51",
         12330 => x"3f",
         12331 => x"08",
         12332 => x"0c",
         12333 => x"04",
         12334 => x"98",
         12335 => x"80",
         12336 => x"08",
         12337 => x"b9",
         12338 => x"33",
         12339 => x"74",
         12340 => x"81",
         12341 => x"38",
         12342 => x"53",
         12343 => x"81",
         12344 => x"fe",
         12345 => x"84",
         12346 => x"80",
         12347 => x"ff",
         12348 => x"75",
         12349 => x"77",
         12350 => x"38",
         12351 => x"58",
         12352 => x"81",
         12353 => x"34",
         12354 => x"7c",
         12355 => x"38",
         12356 => x"51",
         12357 => x"3f",
         12358 => x"08",
         12359 => x"e4",
         12360 => x"ff",
         12361 => x"84",
         12362 => x"06",
         12363 => x"82",
         12364 => x"39",
         12365 => x"17",
         12366 => x"52",
         12367 => x"51",
         12368 => x"3f",
         12369 => x"b8",
         12370 => x"2e",
         12371 => x"ff",
         12372 => x"b8",
         12373 => x"18",
         12374 => x"08",
         12375 => x"31",
         12376 => x"08",
         12377 => x"a0",
         12378 => x"fe",
         12379 => x"17",
         12380 => x"82",
         12381 => x"06",
         12382 => x"81",
         12383 => x"08",
         12384 => x"05",
         12385 => x"81",
         12386 => x"fe",
         12387 => x"79",
         12388 => x"39",
         12389 => x"78",
         12390 => x"38",
         12391 => x"51",
         12392 => x"3f",
         12393 => x"08",
         12394 => x"e4",
         12395 => x"80",
         12396 => x"b8",
         12397 => x"2e",
         12398 => x"84",
         12399 => x"ff",
         12400 => x"38",
         12401 => x"52",
         12402 => x"fd",
         12403 => x"b8",
         12404 => x"38",
         12405 => x"fe",
         12406 => x"08",
         12407 => x"75",
         12408 => x"b0",
         12409 => x"94",
         12410 => x"17",
         12411 => x"5c",
         12412 => x"34",
         12413 => x"7a",
         12414 => x"38",
         12415 => x"a2",
         12416 => x"fd",
         12417 => x"b8",
         12418 => x"fd",
         12419 => x"56",
         12420 => x"e3",
         12421 => x"53",
         12422 => x"bc",
         12423 => x"3d",
         12424 => x"c0",
         12425 => x"e4",
         12426 => x"b8",
         12427 => x"2e",
         12428 => x"84",
         12429 => x"9f",
         12430 => x"7d",
         12431 => x"93",
         12432 => x"5a",
         12433 => x"3f",
         12434 => x"08",
         12435 => x"e4",
         12436 => x"88",
         12437 => x"e4",
         12438 => x"0d",
         12439 => x"e4",
         12440 => x"09",
         12441 => x"38",
         12442 => x"05",
         12443 => x"2a",
         12444 => x"58",
         12445 => x"ff",
         12446 => x"5f",
         12447 => x"3d",
         12448 => x"ff",
         12449 => x"84",
         12450 => x"75",
         12451 => x"b8",
         12452 => x"38",
         12453 => x"b8",
         12454 => x"2e",
         12455 => x"84",
         12456 => x"ff",
         12457 => x"38",
         12458 => x"38",
         12459 => x"e4",
         12460 => x"33",
         12461 => x"7a",
         12462 => x"fe",
         12463 => x"08",
         12464 => x"56",
         12465 => x"79",
         12466 => x"8a",
         12467 => x"71",
         12468 => x"08",
         12469 => x"7a",
         12470 => x"b8",
         12471 => x"80",
         12472 => x"80",
         12473 => x"05",
         12474 => x"15",
         12475 => x"38",
         12476 => x"17",
         12477 => x"75",
         12478 => x"38",
         12479 => x"1b",
         12480 => x"81",
         12481 => x"fe",
         12482 => x"84",
         12483 => x"81",
         12484 => x"18",
         12485 => x"82",
         12486 => x"39",
         12487 => x"17",
         12488 => x"17",
         12489 => x"18",
         12490 => x"fe",
         12491 => x"81",
         12492 => x"e4",
         12493 => x"84",
         12494 => x"83",
         12495 => x"17",
         12496 => x"08",
         12497 => x"a0",
         12498 => x"fe",
         12499 => x"17",
         12500 => x"82",
         12501 => x"06",
         12502 => x"75",
         12503 => x"08",
         12504 => x"05",
         12505 => x"81",
         12506 => x"fe",
         12507 => x"fe",
         12508 => x"56",
         12509 => x"58",
         12510 => x"27",
         12511 => x"7b",
         12512 => x"27",
         12513 => x"74",
         12514 => x"fe",
         12515 => x"84",
         12516 => x"5a",
         12517 => x"08",
         12518 => x"96",
         12519 => x"e4",
         12520 => x"fd",
         12521 => x"b8",
         12522 => x"2e",
         12523 => x"80",
         12524 => x"76",
         12525 => x"b0",
         12526 => x"e4",
         12527 => x"38",
         12528 => x"fe",
         12529 => x"08",
         12530 => x"77",
         12531 => x"38",
         12532 => x"18",
         12533 => x"33",
         12534 => x"7b",
         12535 => x"79",
         12536 => x"26",
         12537 => x"75",
         12538 => x"0c",
         12539 => x"04",
         12540 => x"55",
         12541 => x"ff",
         12542 => x"56",
         12543 => x"09",
         12544 => x"f0",
         12545 => x"b8",
         12546 => x"a0",
         12547 => x"05",
         12548 => x"16",
         12549 => x"38",
         12550 => x"0b",
         12551 => x"7d",
         12552 => x"80",
         12553 => x"7d",
         12554 => x"ce",
         12555 => x"80",
         12556 => x"a1",
         12557 => x"1a",
         12558 => x"0b",
         12559 => x"34",
         12560 => x"ff",
         12561 => x"56",
         12562 => x"17",
         12563 => x"2a",
         12564 => x"d3",
         12565 => x"33",
         12566 => x"2e",
         12567 => x"7d",
         12568 => x"80",
         12569 => x"1b",
         12570 => x"74",
         12571 => x"56",
         12572 => x"81",
         12573 => x"ff",
         12574 => x"ef",
         12575 => x"ae",
         12576 => x"17",
         12577 => x"71",
         12578 => x"06",
         12579 => x"78",
         12580 => x"34",
         12581 => x"5b",
         12582 => x"17",
         12583 => x"55",
         12584 => x"80",
         12585 => x"5b",
         12586 => x"1c",
         12587 => x"ff",
         12588 => x"84",
         12589 => x"56",
         12590 => x"08",
         12591 => x"69",
         12592 => x"e4",
         12593 => x"34",
         12594 => x"08",
         12595 => x"a1",
         12596 => x"34",
         12597 => x"99",
         12598 => x"6a",
         12599 => x"9a",
         12600 => x"88",
         12601 => x"9b",
         12602 => x"33",
         12603 => x"2e",
         12604 => x"69",
         12605 => x"8b",
         12606 => x"57",
         12607 => x"18",
         12608 => x"fe",
         12609 => x"84",
         12610 => x"56",
         12611 => x"e4",
         12612 => x"0d",
         12613 => x"2a",
         12614 => x"ec",
         12615 => x"88",
         12616 => x"80",
         12617 => x"fe",
         12618 => x"90",
         12619 => x"80",
         12620 => x"7a",
         12621 => x"74",
         12622 => x"34",
         12623 => x"0b",
         12624 => x"b8",
         12625 => x"56",
         12626 => x"7b",
         12627 => x"77",
         12628 => x"77",
         12629 => x"7b",
         12630 => x"69",
         12631 => x"8b",
         12632 => x"57",
         12633 => x"18",
         12634 => x"fe",
         12635 => x"84",
         12636 => x"56",
         12637 => x"d1",
         12638 => x"3d",
         12639 => x"70",
         12640 => x"79",
         12641 => x"38",
         12642 => x"05",
         12643 => x"9f",
         12644 => x"75",
         12645 => x"b8",
         12646 => x"38",
         12647 => x"81",
         12648 => x"53",
         12649 => x"fc",
         12650 => x"3d",
         12651 => x"b4",
         12652 => x"e4",
         12653 => x"b8",
         12654 => x"2e",
         12655 => x"84",
         12656 => x"b1",
         12657 => x"7f",
         12658 => x"b2",
         12659 => x"a5",
         12660 => x"59",
         12661 => x"3f",
         12662 => x"08",
         12663 => x"e4",
         12664 => x"02",
         12665 => x"33",
         12666 => x"5d",
         12667 => x"ce",
         12668 => x"92",
         12669 => x"08",
         12670 => x"75",
         12671 => x"57",
         12672 => x"81",
         12673 => x"ff",
         12674 => x"ef",
         12675 => x"58",
         12676 => x"58",
         12677 => x"70",
         12678 => x"33",
         12679 => x"05",
         12680 => x"15",
         12681 => x"38",
         12682 => x"52",
         12683 => x"9e",
         12684 => x"b8",
         12685 => x"84",
         12686 => x"85",
         12687 => x"a8",
         12688 => x"81",
         12689 => x"0b",
         12690 => x"0c",
         12691 => x"04",
         12692 => x"11",
         12693 => x"06",
         12694 => x"74",
         12695 => x"38",
         12696 => x"81",
         12697 => x"05",
         12698 => x"7a",
         12699 => x"38",
         12700 => x"83",
         12701 => x"08",
         12702 => x"5f",
         12703 => x"70",
         12704 => x"33",
         12705 => x"05",
         12706 => x"9f",
         12707 => x"56",
         12708 => x"89",
         12709 => x"70",
         12710 => x"57",
         12711 => x"17",
         12712 => x"26",
         12713 => x"17",
         12714 => x"06",
         12715 => x"30",
         12716 => x"59",
         12717 => x"2e",
         12718 => x"85",
         12719 => x"be",
         12720 => x"32",
         12721 => x"72",
         12722 => x"7a",
         12723 => x"55",
         12724 => x"95",
         12725 => x"84",
         12726 => x"7b",
         12727 => x"c2",
         12728 => x"7e",
         12729 => x"96",
         12730 => x"24",
         12731 => x"79",
         12732 => x"53",
         12733 => x"fc",
         12734 => x"3d",
         12735 => x"e4",
         12736 => x"e4",
         12737 => x"b8",
         12738 => x"b2",
         12739 => x"39",
         12740 => x"08",
         12741 => x"06",
         12742 => x"77",
         12743 => x"a8",
         12744 => x"e4",
         12745 => x"b8",
         12746 => x"92",
         12747 => x"93",
         12748 => x"02",
         12749 => x"cd",
         12750 => x"5a",
         12751 => x"05",
         12752 => x"70",
         12753 => x"34",
         12754 => x"79",
         12755 => x"80",
         12756 => x"8b",
         12757 => x"18",
         12758 => x"2a",
         12759 => x"56",
         12760 => x"75",
         12761 => x"76",
         12762 => x"7f",
         12763 => x"83",
         12764 => x"18",
         12765 => x"2a",
         12766 => x"5c",
         12767 => x"81",
         12768 => x"3d",
         12769 => x"81",
         12770 => x"9b",
         12771 => x"1a",
         12772 => x"2b",
         12773 => x"41",
         12774 => x"7d",
         12775 => x"e0",
         12776 => x"9c",
         12777 => x"05",
         12778 => x"7d",
         12779 => x"38",
         12780 => x"76",
         12781 => x"19",
         12782 => x"5e",
         12783 => x"82",
         12784 => x"7a",
         12785 => x"17",
         12786 => x"aa",
         12787 => x"33",
         12788 => x"bc",
         12789 => x"75",
         12790 => x"52",
         12791 => x"51",
         12792 => x"3f",
         12793 => x"08",
         12794 => x"38",
         12795 => x"5c",
         12796 => x"0c",
         12797 => x"80",
         12798 => x"56",
         12799 => x"38",
         12800 => x"5a",
         12801 => x"09",
         12802 => x"38",
         12803 => x"ff",
         12804 => x"56",
         12805 => x"18",
         12806 => x"2a",
         12807 => x"f3",
         12808 => x"33",
         12809 => x"2e",
         12810 => x"93",
         12811 => x"2a",
         12812 => x"ec",
         12813 => x"88",
         12814 => x"80",
         12815 => x"7f",
         12816 => x"83",
         12817 => x"08",
         12818 => x"b2",
         12819 => x"5c",
         12820 => x"2e",
         12821 => x"52",
         12822 => x"fb",
         12823 => x"b8",
         12824 => x"84",
         12825 => x"80",
         12826 => x"16",
         12827 => x"08",
         12828 => x"b4",
         12829 => x"2e",
         12830 => x"16",
         12831 => x"5f",
         12832 => x"09",
         12833 => x"a8",
         12834 => x"76",
         12835 => x"52",
         12836 => x"51",
         12837 => x"3f",
         12838 => x"08",
         12839 => x"38",
         12840 => x"58",
         12841 => x"0c",
         12842 => x"aa",
         12843 => x"08",
         12844 => x"34",
         12845 => x"17",
         12846 => x"08",
         12847 => x"38",
         12848 => x"51",
         12849 => x"3f",
         12850 => x"08",
         12851 => x"e4",
         12852 => x"ff",
         12853 => x"56",
         12854 => x"f9",
         12855 => x"56",
         12856 => x"38",
         12857 => x"e5",
         12858 => x"b8",
         12859 => x"b8",
         12860 => x"3d",
         12861 => x"0b",
         12862 => x"0c",
         12863 => x"04",
         12864 => x"94",
         12865 => x"98",
         12866 => x"2b",
         12867 => x"58",
         12868 => x"8d",
         12869 => x"e4",
         12870 => x"fb",
         12871 => x"b8",
         12872 => x"2e",
         12873 => x"75",
         12874 => x"0c",
         12875 => x"04",
         12876 => x"16",
         12877 => x"52",
         12878 => x"51",
         12879 => x"3f",
         12880 => x"b8",
         12881 => x"2e",
         12882 => x"fe",
         12883 => x"b8",
         12884 => x"17",
         12885 => x"08",
         12886 => x"31",
         12887 => x"08",
         12888 => x"a0",
         12889 => x"fe",
         12890 => x"16",
         12891 => x"82",
         12892 => x"06",
         12893 => x"81",
         12894 => x"08",
         12895 => x"05",
         12896 => x"81",
         12897 => x"fe",
         12898 => x"79",
         12899 => x"39",
         12900 => x"17",
         12901 => x"17",
         12902 => x"18",
         12903 => x"fe",
         12904 => x"81",
         12905 => x"e4",
         12906 => x"38",
         12907 => x"08",
         12908 => x"b4",
         12909 => x"18",
         12910 => x"b8",
         12911 => x"55",
         12912 => x"08",
         12913 => x"38",
         12914 => x"5d",
         12915 => x"09",
         12916 => x"81",
         12917 => x"b4",
         12918 => x"18",
         12919 => x"7a",
         12920 => x"33",
         12921 => x"eb",
         12922 => x"fb",
         12923 => x"3d",
         12924 => x"df",
         12925 => x"84",
         12926 => x"05",
         12927 => x"82",
         12928 => x"cc",
         12929 => x"3d",
         12930 => x"d8",
         12931 => x"e4",
         12932 => x"b8",
         12933 => x"2e",
         12934 => x"84",
         12935 => x"96",
         12936 => x"78",
         12937 => x"96",
         12938 => x"51",
         12939 => x"3f",
         12940 => x"08",
         12941 => x"e4",
         12942 => x"02",
         12943 => x"33",
         12944 => x"54",
         12945 => x"d2",
         12946 => x"06",
         12947 => x"8b",
         12948 => x"06",
         12949 => x"07",
         12950 => x"55",
         12951 => x"34",
         12952 => x"0b",
         12953 => x"78",
         12954 => x"9a",
         12955 => x"e4",
         12956 => x"e4",
         12957 => x"0d",
         12958 => x"0d",
         12959 => x"53",
         12960 => x"05",
         12961 => x"51",
         12962 => x"3f",
         12963 => x"08",
         12964 => x"e4",
         12965 => x"8a",
         12966 => x"b8",
         12967 => x"3d",
         12968 => x"5a",
         12969 => x"3d",
         12970 => x"ff",
         12971 => x"84",
         12972 => x"55",
         12973 => x"08",
         12974 => x"80",
         12975 => x"81",
         12976 => x"86",
         12977 => x"38",
         12978 => x"22",
         12979 => x"71",
         12980 => x"59",
         12981 => x"96",
         12982 => x"88",
         12983 => x"97",
         12984 => x"90",
         12985 => x"98",
         12986 => x"98",
         12987 => x"99",
         12988 => x"57",
         12989 => x"18",
         12990 => x"fe",
         12991 => x"84",
         12992 => x"84",
         12993 => x"96",
         12994 => x"e8",
         12995 => x"6d",
         12996 => x"53",
         12997 => x"05",
         12998 => x"51",
         12999 => x"3f",
         13000 => x"08",
         13001 => x"08",
         13002 => x"b8",
         13003 => x"80",
         13004 => x"57",
         13005 => x"8b",
         13006 => x"76",
         13007 => x"78",
         13008 => x"76",
         13009 => x"07",
         13010 => x"5b",
         13011 => x"81",
         13012 => x"70",
         13013 => x"58",
         13014 => x"81",
         13015 => x"a4",
         13016 => x"56",
         13017 => x"16",
         13018 => x"82",
         13019 => x"16",
         13020 => x"55",
         13021 => x"09",
         13022 => x"98",
         13023 => x"76",
         13024 => x"52",
         13025 => x"51",
         13026 => x"3f",
         13027 => x"08",
         13028 => x"38",
         13029 => x"59",
         13030 => x"0c",
         13031 => x"bd",
         13032 => x"33",
         13033 => x"c3",
         13034 => x"2e",
         13035 => x"e4",
         13036 => x"2e",
         13037 => x"56",
         13038 => x"05",
         13039 => x"82",
         13040 => x"90",
         13041 => x"2b",
         13042 => x"33",
         13043 => x"88",
         13044 => x"71",
         13045 => x"5f",
         13046 => x"59",
         13047 => x"b8",
         13048 => x"3d",
         13049 => x"5e",
         13050 => x"52",
         13051 => x"52",
         13052 => x"8b",
         13053 => x"e4",
         13054 => x"b8",
         13055 => x"2e",
         13056 => x"76",
         13057 => x"81",
         13058 => x"38",
         13059 => x"80",
         13060 => x"39",
         13061 => x"16",
         13062 => x"16",
         13063 => x"17",
         13064 => x"fe",
         13065 => x"77",
         13066 => x"e4",
         13067 => x"09",
         13068 => x"e8",
         13069 => x"e4",
         13070 => x"34",
         13071 => x"a8",
         13072 => x"84",
         13073 => x"5a",
         13074 => x"17",
         13075 => x"ad",
         13076 => x"33",
         13077 => x"2e",
         13078 => x"fe",
         13079 => x"54",
         13080 => x"a0",
         13081 => x"53",
         13082 => x"16",
         13083 => x"db",
         13084 => x"59",
         13085 => x"53",
         13086 => x"81",
         13087 => x"fe",
         13088 => x"84",
         13089 => x"80",
         13090 => x"38",
         13091 => x"75",
         13092 => x"fe",
         13093 => x"84",
         13094 => x"57",
         13095 => x"08",
         13096 => x"84",
         13097 => x"84",
         13098 => x"66",
         13099 => x"79",
         13100 => x"7c",
         13101 => x"56",
         13102 => x"34",
         13103 => x"8a",
         13104 => x"38",
         13105 => x"57",
         13106 => x"34",
         13107 => x"fc",
         13108 => x"18",
         13109 => x"33",
         13110 => x"79",
         13111 => x"38",
         13112 => x"79",
         13113 => x"39",
         13114 => x"82",
         13115 => x"ff",
         13116 => x"a2",
         13117 => x"9c",
         13118 => x"b8",
         13119 => x"84",
         13120 => x"82",
         13121 => x"3d",
         13122 => x"57",
         13123 => x"70",
         13124 => x"34",
         13125 => x"74",
         13126 => x"a3",
         13127 => x"33",
         13128 => x"06",
         13129 => x"5a",
         13130 => x"81",
         13131 => x"3d",
         13132 => x"5c",
         13133 => x"06",
         13134 => x"55",
         13135 => x"38",
         13136 => x"74",
         13137 => x"26",
         13138 => x"74",
         13139 => x"3f",
         13140 => x"84",
         13141 => x"51",
         13142 => x"84",
         13143 => x"83",
         13144 => x"57",
         13145 => x"81",
         13146 => x"e5",
         13147 => x"e5",
         13148 => x"81",
         13149 => x"56",
         13150 => x"2e",
         13151 => x"74",
         13152 => x"2e",
         13153 => x"18",
         13154 => x"81",
         13155 => x"57",
         13156 => x"2e",
         13157 => x"77",
         13158 => x"06",
         13159 => x"81",
         13160 => x"78",
         13161 => x"81",
         13162 => x"81",
         13163 => x"89",
         13164 => x"38",
         13165 => x"27",
         13166 => x"88",
         13167 => x"7b",
         13168 => x"5d",
         13169 => x"5a",
         13170 => x"81",
         13171 => x"81",
         13172 => x"08",
         13173 => x"81",
         13174 => x"58",
         13175 => x"9f",
         13176 => x"38",
         13177 => x"57",
         13178 => x"81",
         13179 => x"38",
         13180 => x"99",
         13181 => x"05",
         13182 => x"70",
         13183 => x"7a",
         13184 => x"81",
         13185 => x"ff",
         13186 => x"ed",
         13187 => x"80",
         13188 => x"95",
         13189 => x"56",
         13190 => x"3f",
         13191 => x"08",
         13192 => x"e4",
         13193 => x"b4",
         13194 => x"75",
         13195 => x"0c",
         13196 => x"04",
         13197 => x"74",
         13198 => x"3f",
         13199 => x"08",
         13200 => x"06",
         13201 => x"f8",
         13202 => x"75",
         13203 => x"0c",
         13204 => x"04",
         13205 => x"33",
         13206 => x"39",
         13207 => x"51",
         13208 => x"3f",
         13209 => x"08",
         13210 => x"e4",
         13211 => x"38",
         13212 => x"82",
         13213 => x"6c",
         13214 => x"55",
         13215 => x"05",
         13216 => x"70",
         13217 => x"34",
         13218 => x"74",
         13219 => x"5d",
         13220 => x"1e",
         13221 => x"fe",
         13222 => x"84",
         13223 => x"55",
         13224 => x"87",
         13225 => x"27",
         13226 => x"86",
         13227 => x"39",
         13228 => x"08",
         13229 => x"81",
         13230 => x"38",
         13231 => x"75",
         13232 => x"38",
         13233 => x"53",
         13234 => x"fe",
         13235 => x"84",
         13236 => x"57",
         13237 => x"08",
         13238 => x"81",
         13239 => x"38",
         13240 => x"08",
         13241 => x"5a",
         13242 => x"57",
         13243 => x"18",
         13244 => x"b2",
         13245 => x"33",
         13246 => x"2e",
         13247 => x"81",
         13248 => x"54",
         13249 => x"18",
         13250 => x"33",
         13251 => x"c4",
         13252 => x"e4",
         13253 => x"85",
         13254 => x"81",
         13255 => x"19",
         13256 => x"78",
         13257 => x"9c",
         13258 => x"33",
         13259 => x"74",
         13260 => x"81",
         13261 => x"30",
         13262 => x"78",
         13263 => x"74",
         13264 => x"d7",
         13265 => x"5a",
         13266 => x"a5",
         13267 => x"75",
         13268 => x"a1",
         13269 => x"e4",
         13270 => x"b8",
         13271 => x"2e",
         13272 => x"87",
         13273 => x"2e",
         13274 => x"76",
         13275 => x"b9",
         13276 => x"57",
         13277 => x"70",
         13278 => x"34",
         13279 => x"74",
         13280 => x"56",
         13281 => x"17",
         13282 => x"7e",
         13283 => x"76",
         13284 => x"58",
         13285 => x"81",
         13286 => x"ff",
         13287 => x"80",
         13288 => x"38",
         13289 => x"05",
         13290 => x"70",
         13291 => x"34",
         13292 => x"74",
         13293 => x"d6",
         13294 => x"e5",
         13295 => x"5d",
         13296 => x"1e",
         13297 => x"fe",
         13298 => x"84",
         13299 => x"55",
         13300 => x"81",
         13301 => x"39",
         13302 => x"18",
         13303 => x"52",
         13304 => x"51",
         13305 => x"3f",
         13306 => x"08",
         13307 => x"81",
         13308 => x"38",
         13309 => x"08",
         13310 => x"b4",
         13311 => x"19",
         13312 => x"7b",
         13313 => x"27",
         13314 => x"18",
         13315 => x"82",
         13316 => x"84",
         13317 => x"59",
         13318 => x"74",
         13319 => x"75",
         13320 => x"d1",
         13321 => x"e4",
         13322 => x"b8",
         13323 => x"2e",
         13324 => x"fe",
         13325 => x"70",
         13326 => x"80",
         13327 => x"38",
         13328 => x"81",
         13329 => x"08",
         13330 => x"05",
         13331 => x"81",
         13332 => x"fe",
         13333 => x"fd",
         13334 => x"3d",
         13335 => x"02",
         13336 => x"cb",
         13337 => x"5b",
         13338 => x"76",
         13339 => x"38",
         13340 => x"74",
         13341 => x"38",
         13342 => x"73",
         13343 => x"38",
         13344 => x"84",
         13345 => x"59",
         13346 => x"81",
         13347 => x"54",
         13348 => x"81",
         13349 => x"17",
         13350 => x"81",
         13351 => x"80",
         13352 => x"38",
         13353 => x"81",
         13354 => x"17",
         13355 => x"2a",
         13356 => x"5d",
         13357 => x"81",
         13358 => x"8a",
         13359 => x"89",
         13360 => x"7c",
         13361 => x"59",
         13362 => x"3f",
         13363 => x"06",
         13364 => x"72",
         13365 => x"84",
         13366 => x"05",
         13367 => x"79",
         13368 => x"55",
         13369 => x"27",
         13370 => x"19",
         13371 => x"83",
         13372 => x"77",
         13373 => x"80",
         13374 => x"76",
         13375 => x"87",
         13376 => x"7f",
         13377 => x"14",
         13378 => x"83",
         13379 => x"84",
         13380 => x"81",
         13381 => x"38",
         13382 => x"08",
         13383 => x"d8",
         13384 => x"e4",
         13385 => x"38",
         13386 => x"78",
         13387 => x"38",
         13388 => x"09",
         13389 => x"38",
         13390 => x"54",
         13391 => x"e4",
         13392 => x"0d",
         13393 => x"84",
         13394 => x"90",
         13395 => x"81",
         13396 => x"fe",
         13397 => x"84",
         13398 => x"81",
         13399 => x"fe",
         13400 => x"77",
         13401 => x"fe",
         13402 => x"80",
         13403 => x"38",
         13404 => x"58",
         13405 => x"ab",
         13406 => x"54",
         13407 => x"80",
         13408 => x"53",
         13409 => x"51",
         13410 => x"3f",
         13411 => x"08",
         13412 => x"e4",
         13413 => x"38",
         13414 => x"ff",
         13415 => x"5e",
         13416 => x"7e",
         13417 => x"0c",
         13418 => x"2e",
         13419 => x"7a",
         13420 => x"79",
         13421 => x"90",
         13422 => x"c0",
         13423 => x"90",
         13424 => x"15",
         13425 => x"94",
         13426 => x"5a",
         13427 => x"fe",
         13428 => x"7d",
         13429 => x"0c",
         13430 => x"81",
         13431 => x"84",
         13432 => x"54",
         13433 => x"ff",
         13434 => x"39",
         13435 => x"59",
         13436 => x"82",
         13437 => x"39",
         13438 => x"c0",
         13439 => x"5e",
         13440 => x"84",
         13441 => x"e3",
         13442 => x"3d",
         13443 => x"08",
         13444 => x"81",
         13445 => x"44",
         13446 => x"0b",
         13447 => x"70",
         13448 => x"79",
         13449 => x"8a",
         13450 => x"81",
         13451 => x"70",
         13452 => x"56",
         13453 => x"85",
         13454 => x"ed",
         13455 => x"2e",
         13456 => x"84",
         13457 => x"56",
         13458 => x"84",
         13459 => x"10",
         13460 => x"ac",
         13461 => x"56",
         13462 => x"2e",
         13463 => x"75",
         13464 => x"84",
         13465 => x"33",
         13466 => x"12",
         13467 => x"5d",
         13468 => x"51",
         13469 => x"3f",
         13470 => x"08",
         13471 => x"70",
         13472 => x"56",
         13473 => x"84",
         13474 => x"82",
         13475 => x"40",
         13476 => x"84",
         13477 => x"3d",
         13478 => x"83",
         13479 => x"fe",
         13480 => x"84",
         13481 => x"84",
         13482 => x"55",
         13483 => x"84",
         13484 => x"82",
         13485 => x"84",
         13486 => x"15",
         13487 => x"74",
         13488 => x"7e",
         13489 => x"38",
         13490 => x"26",
         13491 => x"7e",
         13492 => x"26",
         13493 => x"ff",
         13494 => x"55",
         13495 => x"38",
         13496 => x"a6",
         13497 => x"2a",
         13498 => x"77",
         13499 => x"5b",
         13500 => x"85",
         13501 => x"30",
         13502 => x"77",
         13503 => x"91",
         13504 => x"b0",
         13505 => x"2e",
         13506 => x"81",
         13507 => x"60",
         13508 => x"fe",
         13509 => x"81",
         13510 => x"e4",
         13511 => x"38",
         13512 => x"05",
         13513 => x"fe",
         13514 => x"88",
         13515 => x"56",
         13516 => x"82",
         13517 => x"09",
         13518 => x"f8",
         13519 => x"29",
         13520 => x"b2",
         13521 => x"58",
         13522 => x"82",
         13523 => x"b6",
         13524 => x"33",
         13525 => x"71",
         13526 => x"88",
         13527 => x"14",
         13528 => x"07",
         13529 => x"33",
         13530 => x"ba",
         13531 => x"33",
         13532 => x"71",
         13533 => x"88",
         13534 => x"14",
         13535 => x"07",
         13536 => x"33",
         13537 => x"a2",
         13538 => x"a3",
         13539 => x"3d",
         13540 => x"54",
         13541 => x"41",
         13542 => x"4d",
         13543 => x"ff",
         13544 => x"90",
         13545 => x"7a",
         13546 => x"82",
         13547 => x"81",
         13548 => x"06",
         13549 => x"80",
         13550 => x"38",
         13551 => x"45",
         13552 => x"89",
         13553 => x"06",
         13554 => x"f4",
         13555 => x"70",
         13556 => x"43",
         13557 => x"83",
         13558 => x"38",
         13559 => x"78",
         13560 => x"81",
         13561 => x"88",
         13562 => x"74",
         13563 => x"38",
         13564 => x"98",
         13565 => x"88",
         13566 => x"82",
         13567 => x"57",
         13568 => x"80",
         13569 => x"76",
         13570 => x"38",
         13571 => x"51",
         13572 => x"3f",
         13573 => x"08",
         13574 => x"55",
         13575 => x"08",
         13576 => x"96",
         13577 => x"84",
         13578 => x"10",
         13579 => x"08",
         13580 => x"72",
         13581 => x"57",
         13582 => x"ff",
         13583 => x"5d",
         13584 => x"47",
         13585 => x"11",
         13586 => x"11",
         13587 => x"6b",
         13588 => x"58",
         13589 => x"62",
         13590 => x"b8",
         13591 => x"5d",
         13592 => x"16",
         13593 => x"56",
         13594 => x"26",
         13595 => x"78",
         13596 => x"31",
         13597 => x"68",
         13598 => x"fd",
         13599 => x"84",
         13600 => x"40",
         13601 => x"89",
         13602 => x"82",
         13603 => x"06",
         13604 => x"83",
         13605 => x"84",
         13606 => x"27",
         13607 => x"7a",
         13608 => x"77",
         13609 => x"80",
         13610 => x"ef",
         13611 => x"fe",
         13612 => x"57",
         13613 => x"e4",
         13614 => x"0d",
         13615 => x"0c",
         13616 => x"fb",
         13617 => x"0b",
         13618 => x"0c",
         13619 => x"84",
         13620 => x"04",
         13621 => x"11",
         13622 => x"06",
         13623 => x"74",
         13624 => x"38",
         13625 => x"81",
         13626 => x"05",
         13627 => x"7a",
         13628 => x"38",
         13629 => x"e4",
         13630 => x"7d",
         13631 => x"5b",
         13632 => x"05",
         13633 => x"70",
         13634 => x"33",
         13635 => x"45",
         13636 => x"99",
         13637 => x"e0",
         13638 => x"ff",
         13639 => x"ff",
         13640 => x"64",
         13641 => x"38",
         13642 => x"81",
         13643 => x"46",
         13644 => x"9f",
         13645 => x"76",
         13646 => x"81",
         13647 => x"78",
         13648 => x"75",
         13649 => x"30",
         13650 => x"9f",
         13651 => x"5d",
         13652 => x"80",
         13653 => x"38",
         13654 => x"1f",
         13655 => x"7c",
         13656 => x"38",
         13657 => x"e0",
         13658 => x"f8",
         13659 => x"52",
         13660 => x"ca",
         13661 => x"57",
         13662 => x"08",
         13663 => x"61",
         13664 => x"06",
         13665 => x"08",
         13666 => x"83",
         13667 => x"6c",
         13668 => x"7e",
         13669 => x"9c",
         13670 => x"31",
         13671 => x"39",
         13672 => x"d2",
         13673 => x"24",
         13674 => x"7b",
         13675 => x"0c",
         13676 => x"39",
         13677 => x"48",
         13678 => x"80",
         13679 => x"38",
         13680 => x"30",
         13681 => x"fc",
         13682 => x"b8",
         13683 => x"f5",
         13684 => x"7a",
         13685 => x"18",
         13686 => x"7b",
         13687 => x"38",
         13688 => x"84",
         13689 => x"9f",
         13690 => x"b8",
         13691 => x"80",
         13692 => x"2e",
         13693 => x"9f",
         13694 => x"8b",
         13695 => x"06",
         13696 => x"7a",
         13697 => x"84",
         13698 => x"55",
         13699 => x"81",
         13700 => x"ff",
         13701 => x"f4",
         13702 => x"83",
         13703 => x"57",
         13704 => x"81",
         13705 => x"76",
         13706 => x"58",
         13707 => x"55",
         13708 => x"60",
         13709 => x"74",
         13710 => x"61",
         13711 => x"77",
         13712 => x"34",
         13713 => x"ff",
         13714 => x"61",
         13715 => x"6a",
         13716 => x"7b",
         13717 => x"34",
         13718 => x"05",
         13719 => x"32",
         13720 => x"48",
         13721 => x"05",
         13722 => x"2a",
         13723 => x"68",
         13724 => x"34",
         13725 => x"83",
         13726 => x"86",
         13727 => x"83",
         13728 => x"55",
         13729 => x"05",
         13730 => x"2a",
         13731 => x"94",
         13732 => x"61",
         13733 => x"bf",
         13734 => x"34",
         13735 => x"05",
         13736 => x"9a",
         13737 => x"61",
         13738 => x"7e",
         13739 => x"34",
         13740 => x"48",
         13741 => x"05",
         13742 => x"2a",
         13743 => x"9e",
         13744 => x"98",
         13745 => x"f0",
         13746 => x"f0",
         13747 => x"05",
         13748 => x"2e",
         13749 => x"80",
         13750 => x"34",
         13751 => x"05",
         13752 => x"a9",
         13753 => x"cc",
         13754 => x"34",
         13755 => x"ff",
         13756 => x"61",
         13757 => x"74",
         13758 => x"6a",
         13759 => x"34",
         13760 => x"a4",
         13761 => x"61",
         13762 => x"93",
         13763 => x"83",
         13764 => x"57",
         13765 => x"81",
         13766 => x"76",
         13767 => x"58",
         13768 => x"55",
         13769 => x"60",
         13770 => x"49",
         13771 => x"34",
         13772 => x"05",
         13773 => x"6b",
         13774 => x"7e",
         13775 => x"79",
         13776 => x"8f",
         13777 => x"84",
         13778 => x"fa",
         13779 => x"17",
         13780 => x"2e",
         13781 => x"69",
         13782 => x"80",
         13783 => x"05",
         13784 => x"15",
         13785 => x"38",
         13786 => x"5b",
         13787 => x"86",
         13788 => x"ff",
         13789 => x"62",
         13790 => x"38",
         13791 => x"61",
         13792 => x"2a",
         13793 => x"74",
         13794 => x"05",
         13795 => x"90",
         13796 => x"64",
         13797 => x"46",
         13798 => x"2a",
         13799 => x"34",
         13800 => x"59",
         13801 => x"83",
         13802 => x"78",
         13803 => x"60",
         13804 => x"fe",
         13805 => x"84",
         13806 => x"85",
         13807 => x"80",
         13808 => x"80",
         13809 => x"05",
         13810 => x"15",
         13811 => x"38",
         13812 => x"7a",
         13813 => x"76",
         13814 => x"81",
         13815 => x"80",
         13816 => x"38",
         13817 => x"83",
         13818 => x"66",
         13819 => x"75",
         13820 => x"38",
         13821 => x"54",
         13822 => x"52",
         13823 => x"c4",
         13824 => x"b8",
         13825 => x"9b",
         13826 => x"76",
         13827 => x"5b",
         13828 => x"8c",
         13829 => x"2e",
         13830 => x"58",
         13831 => x"ff",
         13832 => x"84",
         13833 => x"2e",
         13834 => x"58",
         13835 => x"38",
         13836 => x"81",
         13837 => x"81",
         13838 => x"80",
         13839 => x"80",
         13840 => x"05",
         13841 => x"19",
         13842 => x"38",
         13843 => x"34",
         13844 => x"34",
         13845 => x"05",
         13846 => x"34",
         13847 => x"05",
         13848 => x"82",
         13849 => x"67",
         13850 => x"77",
         13851 => x"34",
         13852 => x"fd",
         13853 => x"1f",
         13854 => x"ab",
         13855 => x"85",
         13856 => x"b8",
         13857 => x"2a",
         13858 => x"76",
         13859 => x"34",
         13860 => x"08",
         13861 => x"34",
         13862 => x"c6",
         13863 => x"61",
         13864 => x"34",
         13865 => x"c8",
         13866 => x"b8",
         13867 => x"83",
         13868 => x"62",
         13869 => x"05",
         13870 => x"2a",
         13871 => x"83",
         13872 => x"62",
         13873 => x"77",
         13874 => x"05",
         13875 => x"2a",
         13876 => x"83",
         13877 => x"81",
         13878 => x"60",
         13879 => x"fe",
         13880 => x"81",
         13881 => x"e4",
         13882 => x"38",
         13883 => x"52",
         13884 => x"c3",
         13885 => x"57",
         13886 => x"08",
         13887 => x"84",
         13888 => x"84",
         13889 => x"9f",
         13890 => x"b8",
         13891 => x"62",
         13892 => x"39",
         13893 => x"16",
         13894 => x"c4",
         13895 => x"38",
         13896 => x"57",
         13897 => x"e6",
         13898 => x"58",
         13899 => x"9d",
         13900 => x"26",
         13901 => x"e6",
         13902 => x"10",
         13903 => x"22",
         13904 => x"74",
         13905 => x"38",
         13906 => x"ee",
         13907 => x"78",
         13908 => x"d3",
         13909 => x"e4",
         13910 => x"84",
         13911 => x"89",
         13912 => x"a0",
         13913 => x"84",
         13914 => x"fc",
         13915 => x"58",
         13916 => x"f0",
         13917 => x"f5",
         13918 => x"57",
         13919 => x"84",
         13920 => x"83",
         13921 => x"f8",
         13922 => x"f8",
         13923 => x"81",
         13924 => x"f4",
         13925 => x"57",
         13926 => x"68",
         13927 => x"63",
         13928 => x"af",
         13929 => x"f4",
         13930 => x"61",
         13931 => x"75",
         13932 => x"68",
         13933 => x"34",
         13934 => x"5b",
         13935 => x"05",
         13936 => x"2a",
         13937 => x"a3",
         13938 => x"c6",
         13939 => x"80",
         13940 => x"80",
         13941 => x"05",
         13942 => x"80",
         13943 => x"80",
         13944 => x"c6",
         13945 => x"61",
         13946 => x"7c",
         13947 => x"7b",
         13948 => x"34",
         13949 => x"59",
         13950 => x"05",
         13951 => x"2a",
         13952 => x"a7",
         13953 => x"61",
         13954 => x"80",
         13955 => x"34",
         13956 => x"05",
         13957 => x"af",
         13958 => x"61",
         13959 => x"80",
         13960 => x"34",
         13961 => x"05",
         13962 => x"b3",
         13963 => x"80",
         13964 => x"05",
         13965 => x"80",
         13966 => x"93",
         13967 => x"05",
         13968 => x"59",
         13969 => x"70",
         13970 => x"33",
         13971 => x"05",
         13972 => x"15",
         13973 => x"2e",
         13974 => x"76",
         13975 => x"58",
         13976 => x"81",
         13977 => x"ff",
         13978 => x"da",
         13979 => x"39",
         13980 => x"53",
         13981 => x"51",
         13982 => x"3f",
         13983 => x"b8",
         13984 => x"b0",
         13985 => x"29",
         13986 => x"77",
         13987 => x"05",
         13988 => x"84",
         13989 => x"53",
         13990 => x"51",
         13991 => x"3f",
         13992 => x"81",
         13993 => x"e4",
         13994 => x"0d",
         13995 => x"0c",
         13996 => x"34",
         13997 => x"6a",
         13998 => x"4c",
         13999 => x"70",
         14000 => x"34",
         14001 => x"ff",
         14002 => x"34",
         14003 => x"05",
         14004 => x"86",
         14005 => x"61",
         14006 => x"ff",
         14007 => x"34",
         14008 => x"05",
         14009 => x"8a",
         14010 => x"65",
         14011 => x"f9",
         14012 => x"54",
         14013 => x"60",
         14014 => x"fe",
         14015 => x"84",
         14016 => x"57",
         14017 => x"81",
         14018 => x"ff",
         14019 => x"f4",
         14020 => x"80",
         14021 => x"81",
         14022 => x"7b",
         14023 => x"75",
         14024 => x"57",
         14025 => x"75",
         14026 => x"57",
         14027 => x"75",
         14028 => x"61",
         14029 => x"34",
         14030 => x"83",
         14031 => x"80",
         14032 => x"e6",
         14033 => x"e1",
         14034 => x"05",
         14035 => x"05",
         14036 => x"83",
         14037 => x"7a",
         14038 => x"78",
         14039 => x"05",
         14040 => x"2a",
         14041 => x"83",
         14042 => x"7a",
         14043 => x"7f",
         14044 => x"05",
         14045 => x"83",
         14046 => x"76",
         14047 => x"05",
         14048 => x"83",
         14049 => x"76",
         14050 => x"05",
         14051 => x"69",
         14052 => x"6b",
         14053 => x"87",
         14054 => x"52",
         14055 => x"bd",
         14056 => x"54",
         14057 => x"60",
         14058 => x"fe",
         14059 => x"69",
         14060 => x"f7",
         14061 => x"3d",
         14062 => x"5b",
         14063 => x"61",
         14064 => x"57",
         14065 => x"25",
         14066 => x"3d",
         14067 => x"f8",
         14068 => x"53",
         14069 => x"51",
         14070 => x"3f",
         14071 => x"09",
         14072 => x"38",
         14073 => x"55",
         14074 => x"90",
         14075 => x"70",
         14076 => x"34",
         14077 => x"74",
         14078 => x"38",
         14079 => x"cd",
         14080 => x"34",
         14081 => x"83",
         14082 => x"74",
         14083 => x"0c",
         14084 => x"04",
         14085 => x"7b",
         14086 => x"b3",
         14087 => x"57",
         14088 => x"80",
         14089 => x"17",
         14090 => x"76",
         14091 => x"88",
         14092 => x"17",
         14093 => x"59",
         14094 => x"81",
         14095 => x"bb",
         14096 => x"74",
         14097 => x"81",
         14098 => x"0c",
         14099 => x"04",
         14100 => x"05",
         14101 => x"8c",
         14102 => x"08",
         14103 => x"d1",
         14104 => x"32",
         14105 => x"72",
         14106 => x"70",
         14107 => x"0c",
         14108 => x"1b",
         14109 => x"56",
         14110 => x"52",
         14111 => x"94",
         14112 => x"39",
         14113 => x"02",
         14114 => x"33",
         14115 => x"58",
         14116 => x"57",
         14117 => x"70",
         14118 => x"34",
         14119 => x"74",
         14120 => x"3d",
         14121 => x"77",
         14122 => x"f7",
         14123 => x"80",
         14124 => x"c0",
         14125 => x"17",
         14126 => x"59",
         14127 => x"81",
         14128 => x"bb",
         14129 => x"74",
         14130 => x"81",
         14131 => x"0c",
         14132 => x"75",
         14133 => x"9f",
         14134 => x"11",
         14135 => x"c0",
         14136 => x"08",
         14137 => x"c9",
         14138 => x"e4",
         14139 => x"7c",
         14140 => x"38",
         14141 => x"b8",
         14142 => x"3d",
         14143 => x"3d",
         14144 => x"55",
         14145 => x"05",
         14146 => x"51",
         14147 => x"3f",
         14148 => x"70",
         14149 => x"07",
         14150 => x"30",
         14151 => x"56",
         14152 => x"8d",
         14153 => x"fd",
         14154 => x"81",
         14155 => x"b8",
         14156 => x"3d",
         14157 => x"3d",
         14158 => x"84",
         14159 => x"22",
         14160 => x"52",
         14161 => x"26",
         14162 => x"83",
         14163 => x"52",
         14164 => x"e4",
         14165 => x"0d",
         14166 => x"ff",
         14167 => x"70",
         14168 => x"09",
         14169 => x"38",
         14170 => x"e4",
         14171 => x"a8",
         14172 => x"71",
         14173 => x"81",
         14174 => x"ff",
         14175 => x"54",
         14176 => x"26",
         14177 => x"10",
         14178 => x"05",
         14179 => x"51",
         14180 => x"80",
         14181 => x"ff",
         14182 => x"e4",
         14183 => x"3d",
         14184 => x"3d",
         14185 => x"05",
         14186 => x"05",
         14187 => x"53",
         14188 => x"70",
         14189 => x"8c",
         14190 => x"72",
         14191 => x"0c",
         14192 => x"04",
         14193 => x"2e",
         14194 => x"ef",
         14195 => x"ff",
         14196 => x"70",
         14197 => x"a8",
         14198 => x"84",
         14199 => x"51",
         14200 => x"04",
         14201 => x"77",
         14202 => x"ff",
         14203 => x"e1",
         14204 => x"ff",
         14205 => x"e8",
         14206 => x"75",
         14207 => x"80",
         14208 => x"70",
         14209 => x"22",
         14210 => x"70",
         14211 => x"7a",
         14212 => x"56",
         14213 => x"b7",
         14214 => x"82",
         14215 => x"72",
         14216 => x"54",
         14217 => x"06",
         14218 => x"54",
         14219 => x"b1",
         14220 => x"38",
         14221 => x"70",
         14222 => x"52",
         14223 => x"30",
         14224 => x"75",
         14225 => x"53",
         14226 => x"80",
         14227 => x"75",
         14228 => x"b8",
         14229 => x"3d",
         14230 => x"ec",
         14231 => x"a2",
         14232 => x"26",
         14233 => x"10",
         14234 => x"d0",
         14235 => x"08",
         14236 => x"16",
         14237 => x"ff",
         14238 => x"75",
         14239 => x"ff",
         14240 => x"83",
         14241 => x"57",
         14242 => x"88",
         14243 => x"ff",
         14244 => x"51",
         14245 => x"16",
         14246 => x"ff",
         14247 => x"db",
         14248 => x"70",
         14249 => x"06",
         14250 => x"39",
         14251 => x"83",
         14252 => x"57",
         14253 => x"f0",
         14254 => x"ff",
         14255 => x"51",
         14256 => x"75",
         14257 => x"06",
         14258 => x"70",
         14259 => x"06",
         14260 => x"ff",
         14261 => x"73",
         14262 => x"05",
         14263 => x"52",
         14264 => x"00",
         14265 => x"ff",
         14266 => x"00",
         14267 => x"ff",
         14268 => x"ff",
         14269 => x"00",
         14270 => x"00",
         14271 => x"00",
         14272 => x"00",
         14273 => x"00",
         14274 => x"00",
         14275 => x"00",
         14276 => x"00",
         14277 => x"00",
         14278 => x"00",
         14279 => x"00",
         14280 => x"00",
         14281 => x"00",
         14282 => x"00",
         14283 => x"00",
         14284 => x"00",
         14285 => x"00",
         14286 => x"00",
         14287 => x"00",
         14288 => x"00",
         14289 => x"00",
         14290 => x"00",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"69",
         14743 => x"00",
         14744 => x"69",
         14745 => x"6c",
         14746 => x"69",
         14747 => x"00",
         14748 => x"6c",
         14749 => x"00",
         14750 => x"65",
         14751 => x"00",
         14752 => x"63",
         14753 => x"72",
         14754 => x"63",
         14755 => x"00",
         14756 => x"64",
         14757 => x"00",
         14758 => x"64",
         14759 => x"00",
         14760 => x"65",
         14761 => x"65",
         14762 => x"65",
         14763 => x"69",
         14764 => x"69",
         14765 => x"66",
         14766 => x"66",
         14767 => x"61",
         14768 => x"00",
         14769 => x"6d",
         14770 => x"65",
         14771 => x"72",
         14772 => x"65",
         14773 => x"00",
         14774 => x"6e",
         14775 => x"00",
         14776 => x"65",
         14777 => x"00",
         14778 => x"6c",
         14779 => x"38",
         14780 => x"62",
         14781 => x"63",
         14782 => x"62",
         14783 => x"63",
         14784 => x"69",
         14785 => x"00",
         14786 => x"64",
         14787 => x"6e",
         14788 => x"77",
         14789 => x"72",
         14790 => x"2e",
         14791 => x"61",
         14792 => x"65",
         14793 => x"73",
         14794 => x"63",
         14795 => x"65",
         14796 => x"00",
         14797 => x"6f",
         14798 => x"61",
         14799 => x"6f",
         14800 => x"20",
         14801 => x"65",
         14802 => x"00",
         14803 => x"6e",
         14804 => x"66",
         14805 => x"65",
         14806 => x"6d",
         14807 => x"72",
         14808 => x"00",
         14809 => x"69",
         14810 => x"69",
         14811 => x"6f",
         14812 => x"64",
         14813 => x"69",
         14814 => x"75",
         14815 => x"6f",
         14816 => x"61",
         14817 => x"6e",
         14818 => x"6e",
         14819 => x"6c",
         14820 => x"00",
         14821 => x"6f",
         14822 => x"74",
         14823 => x"6f",
         14824 => x"64",
         14825 => x"6f",
         14826 => x"6d",
         14827 => x"69",
         14828 => x"20",
         14829 => x"65",
         14830 => x"74",
         14831 => x"66",
         14832 => x"64",
         14833 => x"20",
         14834 => x"6b",
         14835 => x"69",
         14836 => x"6e",
         14837 => x"65",
         14838 => x"6c",
         14839 => x"00",
         14840 => x"72",
         14841 => x"20",
         14842 => x"62",
         14843 => x"69",
         14844 => x"6e",
         14845 => x"69",
         14846 => x"00",
         14847 => x"44",
         14848 => x"20",
         14849 => x"74",
         14850 => x"72",
         14851 => x"63",
         14852 => x"2e",
         14853 => x"69",
         14854 => x"68",
         14855 => x"6c",
         14856 => x"6e",
         14857 => x"69",
         14858 => x"00",
         14859 => x"69",
         14860 => x"61",
         14861 => x"61",
         14862 => x"65",
         14863 => x"74",
         14864 => x"00",
         14865 => x"63",
         14866 => x"73",
         14867 => x"6e",
         14868 => x"2e",
         14869 => x"6e",
         14870 => x"69",
         14871 => x"69",
         14872 => x"61",
         14873 => x"00",
         14874 => x"6f",
         14875 => x"74",
         14876 => x"6f",
         14877 => x"2e",
         14878 => x"6f",
         14879 => x"6c",
         14880 => x"6f",
         14881 => x"2e",
         14882 => x"69",
         14883 => x"6e",
         14884 => x"72",
         14885 => x"79",
         14886 => x"6e",
         14887 => x"6e",
         14888 => x"65",
         14889 => x"72",
         14890 => x"69",
         14891 => x"45",
         14892 => x"72",
         14893 => x"75",
         14894 => x"73",
         14895 => x"00",
         14896 => x"25",
         14897 => x"62",
         14898 => x"73",
         14899 => x"20",
         14900 => x"25",
         14901 => x"62",
         14902 => x"73",
         14903 => x"63",
         14904 => x"00",
         14905 => x"65",
         14906 => x"00",
         14907 => x"30",
         14908 => x"00",
         14909 => x"20",
         14910 => x"30",
         14911 => x"00",
         14912 => x"7c",
         14913 => x"00",
         14914 => x"20",
         14915 => x"30",
         14916 => x"00",
         14917 => x"20",
         14918 => x"20",
         14919 => x"00",
         14920 => x"4f",
         14921 => x"2a",
         14922 => x"20",
         14923 => x"37",
         14924 => x"2f",
         14925 => x"31",
         14926 => x"31",
         14927 => x"00",
         14928 => x"5a",
         14929 => x"20",
         14930 => x"20",
         14931 => x"78",
         14932 => x"73",
         14933 => x"20",
         14934 => x"0a",
         14935 => x"50",
         14936 => x"6e",
         14937 => x"72",
         14938 => x"20",
         14939 => x"64",
         14940 => x"00",
         14941 => x"41",
         14942 => x"20",
         14943 => x"69",
         14944 => x"72",
         14945 => x"74",
         14946 => x"41",
         14947 => x"20",
         14948 => x"69",
         14949 => x"72",
         14950 => x"74",
         14951 => x"41",
         14952 => x"20",
         14953 => x"69",
         14954 => x"72",
         14955 => x"74",
         14956 => x"41",
         14957 => x"20",
         14958 => x"69",
         14959 => x"72",
         14960 => x"74",
         14961 => x"4f",
         14962 => x"20",
         14963 => x"69",
         14964 => x"72",
         14965 => x"74",
         14966 => x"4f",
         14967 => x"20",
         14968 => x"69",
         14969 => x"72",
         14970 => x"74",
         14971 => x"53",
         14972 => x"6e",
         14973 => x"72",
         14974 => x"00",
         14975 => x"69",
         14976 => x"20",
         14977 => x"65",
         14978 => x"70",
         14979 => x"65",
         14980 => x"6e",
         14981 => x"70",
         14982 => x"6d",
         14983 => x"2e",
         14984 => x"6e",
         14985 => x"69",
         14986 => x"74",
         14987 => x"72",
         14988 => x"00",
         14989 => x"75",
         14990 => x"78",
         14991 => x"62",
         14992 => x"00",
         14993 => x"4f",
         14994 => x"70",
         14995 => x"73",
         14996 => x"61",
         14997 => x"64",
         14998 => x"20",
         14999 => x"74",
         15000 => x"69",
         15001 => x"73",
         15002 => x"61",
         15003 => x"30",
         15004 => x"6c",
         15005 => x"65",
         15006 => x"69",
         15007 => x"61",
         15008 => x"6c",
         15009 => x"00",
         15010 => x"20",
         15011 => x"64",
         15012 => x"73",
         15013 => x"3a",
         15014 => x"61",
         15015 => x"6f",
         15016 => x"6e",
         15017 => x"00",
         15018 => x"50",
         15019 => x"69",
         15020 => x"64",
         15021 => x"73",
         15022 => x"2e",
         15023 => x"00",
         15024 => x"6f",
         15025 => x"72",
         15026 => x"6f",
         15027 => x"67",
         15028 => x"00",
         15029 => x"65",
         15030 => x"72",
         15031 => x"67",
         15032 => x"70",
         15033 => x"61",
         15034 => x"6e",
         15035 => x"00",
         15036 => x"61",
         15037 => x"6e",
         15038 => x"6f",
         15039 => x"40",
         15040 => x"38",
         15041 => x"2e",
         15042 => x"00",
         15043 => x"61",
         15044 => x"72",
         15045 => x"72",
         15046 => x"20",
         15047 => x"65",
         15048 => x"64",
         15049 => x"00",
         15050 => x"78",
         15051 => x"74",
         15052 => x"20",
         15053 => x"65",
         15054 => x"25",
         15055 => x"78",
         15056 => x"2e",
         15057 => x"30",
         15058 => x"20",
         15059 => x"6c",
         15060 => x"00",
         15061 => x"30",
         15062 => x"20",
         15063 => x"58",
         15064 => x"6f",
         15065 => x"72",
         15066 => x"2e",
         15067 => x"00",
         15068 => x"30",
         15069 => x"28",
         15070 => x"78",
         15071 => x"25",
         15072 => x"78",
         15073 => x"38",
         15074 => x"00",
         15075 => x"6f",
         15076 => x"6e",
         15077 => x"2e",
         15078 => x"30",
         15079 => x"20",
         15080 => x"58",
         15081 => x"6c",
         15082 => x"69",
         15083 => x"2e",
         15084 => x"00",
         15085 => x"75",
         15086 => x"4d",
         15087 => x"72",
         15088 => x"43",
         15089 => x"6c",
         15090 => x"2e",
         15091 => x"64",
         15092 => x"73",
         15093 => x"00",
         15094 => x"65",
         15095 => x"79",
         15096 => x"68",
         15097 => x"74",
         15098 => x"20",
         15099 => x"6e",
         15100 => x"70",
         15101 => x"65",
         15102 => x"63",
         15103 => x"61",
         15104 => x"00",
         15105 => x"3f",
         15106 => x"64",
         15107 => x"2f",
         15108 => x"25",
         15109 => x"64",
         15110 => x"2e",
         15111 => x"64",
         15112 => x"6f",
         15113 => x"6f",
         15114 => x"67",
         15115 => x"74",
         15116 => x"00",
         15117 => x"0a",
         15118 => x"69",
         15119 => x"20",
         15120 => x"6c",
         15121 => x"6e",
         15122 => x"3a",
         15123 => x"64",
         15124 => x"73",
         15125 => x"3a",
         15126 => x"20",
         15127 => x"50",
         15128 => x"65",
         15129 => x"20",
         15130 => x"74",
         15131 => x"41",
         15132 => x"65",
         15133 => x"3d",
         15134 => x"38",
         15135 => x"00",
         15136 => x"20",
         15137 => x"50",
         15138 => x"65",
         15139 => x"79",
         15140 => x"61",
         15141 => x"41",
         15142 => x"65",
         15143 => x"3d",
         15144 => x"38",
         15145 => x"00",
         15146 => x"20",
         15147 => x"74",
         15148 => x"20",
         15149 => x"72",
         15150 => x"64",
         15151 => x"73",
         15152 => x"20",
         15153 => x"3d",
         15154 => x"38",
         15155 => x"00",
         15156 => x"69",
         15157 => x"00",
         15158 => x"20",
         15159 => x"50",
         15160 => x"64",
         15161 => x"20",
         15162 => x"20",
         15163 => x"20",
         15164 => x"20",
         15165 => x"3d",
         15166 => x"34",
         15167 => x"00",
         15168 => x"20",
         15169 => x"79",
         15170 => x"6d",
         15171 => x"6f",
         15172 => x"46",
         15173 => x"20",
         15174 => x"20",
         15175 => x"3d",
         15176 => x"2e",
         15177 => x"64",
         15178 => x"0a",
         15179 => x"20",
         15180 => x"69",
         15181 => x"6f",
         15182 => x"53",
         15183 => x"4d",
         15184 => x"6f",
         15185 => x"46",
         15186 => x"3d",
         15187 => x"2e",
         15188 => x"64",
         15189 => x"0a",
         15190 => x"20",
         15191 => x"44",
         15192 => x"20",
         15193 => x"63",
         15194 => x"72",
         15195 => x"20",
         15196 => x"20",
         15197 => x"3d",
         15198 => x"2e",
         15199 => x"64",
         15200 => x"0a",
         15201 => x"20",
         15202 => x"50",
         15203 => x"20",
         15204 => x"53",
         15205 => x"20",
         15206 => x"4f",
         15207 => x"00",
         15208 => x"20",
         15209 => x"42",
         15210 => x"43",
         15211 => x"20",
         15212 => x"49",
         15213 => x"4f",
         15214 => x"42",
         15215 => x"00",
         15216 => x"20",
         15217 => x"4e",
         15218 => x"43",
         15219 => x"20",
         15220 => x"61",
         15221 => x"6c",
         15222 => x"30",
         15223 => x"2e",
         15224 => x"20",
         15225 => x"49",
         15226 => x"31",
         15227 => x"20",
         15228 => x"6d",
         15229 => x"20",
         15230 => x"30",
         15231 => x"2e",
         15232 => x"20",
         15233 => x"44",
         15234 => x"52",
         15235 => x"20",
         15236 => x"76",
         15237 => x"73",
         15238 => x"30",
         15239 => x"2e",
         15240 => x"20",
         15241 => x"41",
         15242 => x"20",
         15243 => x"20",
         15244 => x"38",
         15245 => x"30",
         15246 => x"2e",
         15247 => x"20",
         15248 => x"52",
         15249 => x"20",
         15250 => x"20",
         15251 => x"38",
         15252 => x"30",
         15253 => x"2e",
         15254 => x"20",
         15255 => x"4e",
         15256 => x"42",
         15257 => x"20",
         15258 => x"38",
         15259 => x"30",
         15260 => x"2e",
         15261 => x"20",
         15262 => x"44",
         15263 => x"20",
         15264 => x"20",
         15265 => x"38",
         15266 => x"30",
         15267 => x"2e",
         15268 => x"20",
         15269 => x"42",
         15270 => x"52",
         15271 => x"20",
         15272 => x"38",
         15273 => x"30",
         15274 => x"2e",
         15275 => x"28",
         15276 => x"6d",
         15277 => x"43",
         15278 => x"6e",
         15279 => x"29",
         15280 => x"6e",
         15281 => x"77",
         15282 => x"56",
         15283 => x"00",
         15284 => x"6d",
         15285 => x"00",
         15286 => x"65",
         15287 => x"6d",
         15288 => x"6c",
         15289 => x"00",
         15290 => x"56",
         15291 => x"00",
         15292 => x"00",
         15293 => x"00",
         15294 => x"00",
         15295 => x"00",
         15296 => x"00",
         15297 => x"00",
         15298 => x"00",
         15299 => x"00",
         15300 => x"00",
         15301 => x"00",
         15302 => x"00",
         15303 => x"00",
         15304 => x"00",
         15305 => x"00",
         15306 => x"00",
         15307 => x"00",
         15308 => x"00",
         15309 => x"00",
         15310 => x"00",
         15311 => x"00",
         15312 => x"00",
         15313 => x"00",
         15314 => x"00",
         15315 => x"00",
         15316 => x"00",
         15317 => x"00",
         15318 => x"00",
         15319 => x"00",
         15320 => x"00",
         15321 => x"00",
         15322 => x"00",
         15323 => x"00",
         15324 => x"00",
         15325 => x"00",
         15326 => x"00",
         15327 => x"00",
         15328 => x"00",
         15329 => x"00",
         15330 => x"00",
         15331 => x"00",
         15332 => x"00",
         15333 => x"00",
         15334 => x"00",
         15335 => x"00",
         15336 => x"00",
         15337 => x"00",
         15338 => x"00",
         15339 => x"00",
         15340 => x"00",
         15341 => x"00",
         15342 => x"00",
         15343 => x"00",
         15344 => x"00",
         15345 => x"00",
         15346 => x"00",
         15347 => x"00",
         15348 => x"00",
         15349 => x"00",
         15350 => x"00",
         15351 => x"00",
         15352 => x"00",
         15353 => x"00",
         15354 => x"00",
         15355 => x"00",
         15356 => x"00",
         15357 => x"5b",
         15358 => x"5b",
         15359 => x"5b",
         15360 => x"5b",
         15361 => x"5b",
         15362 => x"5b",
         15363 => x"5b",
         15364 => x"30",
         15365 => x"5b",
         15366 => x"5b",
         15367 => x"5b",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"61",
         15380 => x"74",
         15381 => x"65",
         15382 => x"72",
         15383 => x"65",
         15384 => x"73",
         15385 => x"79",
         15386 => x"6c",
         15387 => x"64",
         15388 => x"62",
         15389 => x"67",
         15390 => x"69",
         15391 => x"72",
         15392 => x"69",
         15393 => x"00",
         15394 => x"00",
         15395 => x"30",
         15396 => x"20",
         15397 => x"0a",
         15398 => x"61",
         15399 => x"64",
         15400 => x"20",
         15401 => x"65",
         15402 => x"68",
         15403 => x"69",
         15404 => x"72",
         15405 => x"69",
         15406 => x"74",
         15407 => x"4f",
         15408 => x"00",
         15409 => x"25",
         15410 => x"00",
         15411 => x"5b",
         15412 => x"00",
         15413 => x"5b",
         15414 => x"5b",
         15415 => x"5b",
         15416 => x"5b",
         15417 => x"5b",
         15418 => x"00",
         15419 => x"5b",
         15420 => x"00",
         15421 => x"5b",
         15422 => x"00",
         15423 => x"5b",
         15424 => x"00",
         15425 => x"5b",
         15426 => x"00",
         15427 => x"5b",
         15428 => x"00",
         15429 => x"5b",
         15430 => x"00",
         15431 => x"5b",
         15432 => x"00",
         15433 => x"5b",
         15434 => x"00",
         15435 => x"5b",
         15436 => x"00",
         15437 => x"5b",
         15438 => x"00",
         15439 => x"5b",
         15440 => x"00",
         15441 => x"5b",
         15442 => x"5b",
         15443 => x"00",
         15444 => x"5b",
         15445 => x"00",
         15446 => x"3a",
         15447 => x"25",
         15448 => x"64",
         15449 => x"2c",
         15450 => x"25",
         15451 => x"30",
         15452 => x"00",
         15453 => x"3a",
         15454 => x"25",
         15455 => x"64",
         15456 => x"3a",
         15457 => x"25",
         15458 => x"64",
         15459 => x"64",
         15460 => x"3a",
         15461 => x"00",
         15462 => x"30",
         15463 => x"00",
         15464 => x"63",
         15465 => x"3b",
         15466 => x"00",
         15467 => x"65",
         15468 => x"74",
         15469 => x"72",
         15470 => x"3a",
         15471 => x"70",
         15472 => x"32",
         15473 => x"30",
         15474 => x"00",
         15475 => x"77",
         15476 => x"32",
         15477 => x"30",
         15478 => x"00",
         15479 => x"64",
         15480 => x"32",
         15481 => x"00",
         15482 => x"6f",
         15483 => x"73",
         15484 => x"65",
         15485 => x"65",
         15486 => x"00",
         15487 => x"44",
         15488 => x"2a",
         15489 => x"3f",
         15490 => x"00",
         15491 => x"2c",
         15492 => x"5d",
         15493 => x"41",
         15494 => x"41",
         15495 => x"00",
         15496 => x"fe",
         15497 => x"44",
         15498 => x"2e",
         15499 => x"4f",
         15500 => x"4d",
         15501 => x"20",
         15502 => x"54",
         15503 => x"20",
         15504 => x"4f",
         15505 => x"4d",
         15506 => x"20",
         15507 => x"54",
         15508 => x"20",
         15509 => x"00",
         15510 => x"00",
         15511 => x"00",
         15512 => x"00",
         15513 => x"03",
         15514 => x"0e",
         15515 => x"16",
         15516 => x"00",
         15517 => x"9a",
         15518 => x"41",
         15519 => x"45",
         15520 => x"49",
         15521 => x"92",
         15522 => x"4f",
         15523 => x"99",
         15524 => x"9d",
         15525 => x"49",
         15526 => x"a5",
         15527 => x"a9",
         15528 => x"ad",
         15529 => x"b1",
         15530 => x"b5",
         15531 => x"b9",
         15532 => x"bd",
         15533 => x"c1",
         15534 => x"c5",
         15535 => x"c9",
         15536 => x"cd",
         15537 => x"d1",
         15538 => x"d5",
         15539 => x"d9",
         15540 => x"dd",
         15541 => x"e1",
         15542 => x"e5",
         15543 => x"e9",
         15544 => x"ed",
         15545 => x"f1",
         15546 => x"f5",
         15547 => x"f9",
         15548 => x"fd",
         15549 => x"2e",
         15550 => x"5b",
         15551 => x"22",
         15552 => x"3e",
         15553 => x"00",
         15554 => x"01",
         15555 => x"10",
         15556 => x"00",
         15557 => x"00",
         15558 => x"01",
         15559 => x"04",
         15560 => x"10",
         15561 => x"00",
         15562 => x"c7",
         15563 => x"e9",
         15564 => x"e4",
         15565 => x"e5",
         15566 => x"ea",
         15567 => x"e8",
         15568 => x"ee",
         15569 => x"c4",
         15570 => x"c9",
         15571 => x"c6",
         15572 => x"f6",
         15573 => x"fb",
         15574 => x"ff",
         15575 => x"dc",
         15576 => x"a3",
         15577 => x"a7",
         15578 => x"e1",
         15579 => x"f3",
         15580 => x"f1",
         15581 => x"aa",
         15582 => x"bf",
         15583 => x"ac",
         15584 => x"bc",
         15585 => x"ab",
         15586 => x"91",
         15587 => x"93",
         15588 => x"24",
         15589 => x"62",
         15590 => x"55",
         15591 => x"51",
         15592 => x"5d",
         15593 => x"5b",
         15594 => x"14",
         15595 => x"2c",
         15596 => x"00",
         15597 => x"5e",
         15598 => x"5a",
         15599 => x"69",
         15600 => x"60",
         15601 => x"6c",
         15602 => x"68",
         15603 => x"65",
         15604 => x"58",
         15605 => x"53",
         15606 => x"6a",
         15607 => x"0c",
         15608 => x"84",
         15609 => x"90",
         15610 => x"b1",
         15611 => x"93",
         15612 => x"a3",
         15613 => x"b5",
         15614 => x"a6",
         15615 => x"a9",
         15616 => x"1e",
         15617 => x"b5",
         15618 => x"61",
         15619 => x"65",
         15620 => x"20",
         15621 => x"f7",
         15622 => x"b0",
         15623 => x"b7",
         15624 => x"7f",
         15625 => x"a0",
         15626 => x"61",
         15627 => x"e0",
         15628 => x"f8",
         15629 => x"ff",
         15630 => x"78",
         15631 => x"30",
         15632 => x"06",
         15633 => x"10",
         15634 => x"2e",
         15635 => x"06",
         15636 => x"4d",
         15637 => x"81",
         15638 => x"82",
         15639 => x"84",
         15640 => x"87",
         15641 => x"89",
         15642 => x"8b",
         15643 => x"8d",
         15644 => x"8f",
         15645 => x"91",
         15646 => x"93",
         15647 => x"f6",
         15648 => x"97",
         15649 => x"98",
         15650 => x"9b",
         15651 => x"9d",
         15652 => x"9f",
         15653 => x"a0",
         15654 => x"a2",
         15655 => x"a4",
         15656 => x"a7",
         15657 => x"a9",
         15658 => x"ab",
         15659 => x"ac",
         15660 => x"af",
         15661 => x"b1",
         15662 => x"b3",
         15663 => x"b5",
         15664 => x"b7",
         15665 => x"b8",
         15666 => x"bb",
         15667 => x"bc",
         15668 => x"f7",
         15669 => x"c1",
         15670 => x"c3",
         15671 => x"c5",
         15672 => x"c7",
         15673 => x"c7",
         15674 => x"cb",
         15675 => x"cd",
         15676 => x"dd",
         15677 => x"8e",
         15678 => x"12",
         15679 => x"03",
         15680 => x"f4",
         15681 => x"f8",
         15682 => x"22",
         15683 => x"3a",
         15684 => x"65",
         15685 => x"3b",
         15686 => x"66",
         15687 => x"40",
         15688 => x"41",
         15689 => x"0a",
         15690 => x"40",
         15691 => x"86",
         15692 => x"89",
         15693 => x"58",
         15694 => x"5a",
         15695 => x"5c",
         15696 => x"5e",
         15697 => x"93",
         15698 => x"62",
         15699 => x"64",
         15700 => x"66",
         15701 => x"97",
         15702 => x"6a",
         15703 => x"6c",
         15704 => x"6e",
         15705 => x"70",
         15706 => x"9d",
         15707 => x"74",
         15708 => x"76",
         15709 => x"78",
         15710 => x"7a",
         15711 => x"7c",
         15712 => x"7e",
         15713 => x"a6",
         15714 => x"82",
         15715 => x"84",
         15716 => x"86",
         15717 => x"ae",
         15718 => x"b1",
         15719 => x"45",
         15720 => x"8e",
         15721 => x"90",
         15722 => x"b7",
         15723 => x"03",
         15724 => x"fe",
         15725 => x"ac",
         15726 => x"86",
         15727 => x"89",
         15728 => x"b1",
         15729 => x"c2",
         15730 => x"a3",
         15731 => x"c4",
         15732 => x"cc",
         15733 => x"8c",
         15734 => x"8f",
         15735 => x"18",
         15736 => x"0a",
         15737 => x"f3",
         15738 => x"f5",
         15739 => x"f7",
         15740 => x"f9",
         15741 => x"fa",
         15742 => x"20",
         15743 => x"10",
         15744 => x"22",
         15745 => x"36",
         15746 => x"0e",
         15747 => x"01",
         15748 => x"d0",
         15749 => x"61",
         15750 => x"00",
         15751 => x"7d",
         15752 => x"63",
         15753 => x"96",
         15754 => x"5a",
         15755 => x"08",
         15756 => x"06",
         15757 => x"08",
         15758 => x"08",
         15759 => x"06",
         15760 => x"07",
         15761 => x"52",
         15762 => x"54",
         15763 => x"56",
         15764 => x"60",
         15765 => x"70",
         15766 => x"ba",
         15767 => x"c8",
         15768 => x"ca",
         15769 => x"da",
         15770 => x"f8",
         15771 => x"ea",
         15772 => x"fa",
         15773 => x"80",
         15774 => x"90",
         15775 => x"a0",
         15776 => x"b0",
         15777 => x"b8",
         15778 => x"b2",
         15779 => x"cc",
         15780 => x"c3",
         15781 => x"02",
         15782 => x"02",
         15783 => x"01",
         15784 => x"f3",
         15785 => x"fc",
         15786 => x"01",
         15787 => x"70",
         15788 => x"84",
         15789 => x"83",
         15790 => x"1a",
         15791 => x"2f",
         15792 => x"02",
         15793 => x"06",
         15794 => x"02",
         15795 => x"64",
         15796 => x"26",
         15797 => x"1a",
         15798 => x"00",
         15799 => x"00",
         15800 => x"02",
         15801 => x"00",
         15802 => x"00",
         15803 => x"00",
         15804 => x"04",
         15805 => x"00",
         15806 => x"00",
         15807 => x"00",
         15808 => x"14",
         15809 => x"00",
         15810 => x"00",
         15811 => x"00",
         15812 => x"2b",
         15813 => x"00",
         15814 => x"00",
         15815 => x"00",
         15816 => x"30",
         15817 => x"00",
         15818 => x"00",
         15819 => x"00",
         15820 => x"3c",
         15821 => x"00",
         15822 => x"00",
         15823 => x"00",
         15824 => x"3d",
         15825 => x"00",
         15826 => x"00",
         15827 => x"00",
         15828 => x"3f",
         15829 => x"00",
         15830 => x"00",
         15831 => x"00",
         15832 => x"40",
         15833 => x"00",
         15834 => x"00",
         15835 => x"00",
         15836 => x"41",
         15837 => x"00",
         15838 => x"00",
         15839 => x"00",
         15840 => x"42",
         15841 => x"00",
         15842 => x"00",
         15843 => x"00",
         15844 => x"43",
         15845 => x"00",
         15846 => x"00",
         15847 => x"00",
         15848 => x"50",
         15849 => x"00",
         15850 => x"00",
         15851 => x"00",
         15852 => x"51",
         15853 => x"00",
         15854 => x"00",
         15855 => x"00",
         15856 => x"54",
         15857 => x"00",
         15858 => x"00",
         15859 => x"00",
         15860 => x"55",
         15861 => x"00",
         15862 => x"00",
         15863 => x"00",
         15864 => x"79",
         15865 => x"00",
         15866 => x"00",
         15867 => x"00",
         15868 => x"78",
         15869 => x"00",
         15870 => x"00",
         15871 => x"00",
         15872 => x"82",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"83",
         15877 => x"00",
         15878 => x"00",
         15879 => x"00",
         15880 => x"85",
         15881 => x"00",
         15882 => x"00",
         15883 => x"00",
         15884 => x"87",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"88",
         15889 => x"00",
         15890 => x"00",
         15891 => x"00",
         15892 => x"89",
         15893 => x"00",
         15894 => x"00",
         15895 => x"00",
         15896 => x"8c",
         15897 => x"00",
         15898 => x"00",
         15899 => x"00",
         15900 => x"8d",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"8e",
         15905 => x"00",
         15906 => x"00",
         15907 => x"00",
         15908 => x"8f",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"00",
         15914 => x"00",
         15915 => x"00",
         15916 => x"01",
         15917 => x"00",
         15918 => x"01",
         15919 => x"81",
         15920 => x"00",
         15921 => x"7f",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"00",
         15926 => x"f5",
         15927 => x"f5",
         15928 => x"f5",
         15929 => x"00",
         15930 => x"01",
         15931 => x"01",
         15932 => x"01",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"00",
         15959 => x"00",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"01",
         15965 => x"fc",
         15966 => x"3b",
         15967 => x"7a",
         15968 => x"f0",
         15969 => x"72",
         15970 => x"76",
         15971 => x"6a",
         15972 => x"6e",
         15973 => x"62",
         15974 => x"66",
         15975 => x"32",
         15976 => x"36",
         15977 => x"f3",
         15978 => x"39",
         15979 => x"7f",
         15980 => x"f2",
         15981 => x"f0",
         15982 => x"f0",
         15983 => x"81",
         15984 => x"f0",
         15985 => x"fc",
         15986 => x"3a",
         15987 => x"5a",
         15988 => x"f0",
         15989 => x"52",
         15990 => x"56",
         15991 => x"4a",
         15992 => x"4e",
         15993 => x"42",
         15994 => x"46",
         15995 => x"32",
         15996 => x"36",
         15997 => x"f3",
         15998 => x"39",
         15999 => x"7f",
         16000 => x"f2",
         16001 => x"f0",
         16002 => x"f0",
         16003 => x"81",
         16004 => x"f0",
         16005 => x"fc",
         16006 => x"2b",
         16007 => x"5a",
         16008 => x"f0",
         16009 => x"52",
         16010 => x"56",
         16011 => x"4a",
         16012 => x"4e",
         16013 => x"42",
         16014 => x"46",
         16015 => x"22",
         16016 => x"26",
         16017 => x"7e",
         16018 => x"29",
         16019 => x"e2",
         16020 => x"f8",
         16021 => x"f0",
         16022 => x"f0",
         16023 => x"86",
         16024 => x"f0",
         16025 => x"fe",
         16026 => x"f0",
         16027 => x"1a",
         16028 => x"f0",
         16029 => x"12",
         16030 => x"16",
         16031 => x"0a",
         16032 => x"0e",
         16033 => x"02",
         16034 => x"06",
         16035 => x"f0",
         16036 => x"f0",
         16037 => x"1e",
         16038 => x"1f",
         16039 => x"f0",
         16040 => x"f0",
         16041 => x"f0",
         16042 => x"f0",
         16043 => x"81",
         16044 => x"f0",
         16045 => x"f0",
         16046 => x"b5",
         16047 => x"77",
         16048 => x"f0",
         16049 => x"70",
         16050 => x"a6",
         16051 => x"5d",
         16052 => x"33",
         16053 => x"6e",
         16054 => x"43",
         16055 => x"36",
         16056 => x"1e",
         16057 => x"9f",
         16058 => x"a3",
         16059 => x"c5",
         16060 => x"c4",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"81",
         16064 => x"f0",
         16065 => x"00",
         16066 => x"00",
         16067 => x"00",
         16068 => x"00",
         16069 => x"00",
         16070 => x"00",
         16071 => x"00",
         16072 => x"00",
         16073 => x"00",
         16074 => x"00",
         16075 => x"00",
         16076 => x"00",
         16077 => x"00",
         16078 => x"00",
         16079 => x"00",
         16080 => x"00",
         16081 => x"00",
         16082 => x"00",
         16083 => x"00",
         16084 => x"00",
         16085 => x"00",
         16086 => x"00",
         16087 => x"00",
         16088 => x"00",
         16089 => x"00",
         16090 => x"01",
         16091 => x"00",
         16092 => x"00",
         16093 => x"00",
         16094 => x"00",
         16095 => x"00",
         16096 => x"00",
         16097 => x"00",
         16098 => x"00",
         16099 => x"00",
         16100 => x"00",
         16101 => x"00",
         16102 => x"00",
         16103 => x"00",
         16104 => x"00",
         16105 => x"00",
         16106 => x"00",
         16107 => x"00",
         16108 => x"00",
         16109 => x"00",
         16110 => x"00",
         16111 => x"00",
         16112 => x"00",
         16113 => x"00",
         16114 => x"00",
         16115 => x"00",
         16116 => x"00",
         16117 => x"00",
         16118 => x"00",
         16119 => x"00",
         16120 => x"00",
         16121 => x"00",
         16122 => x"00",
         16123 => x"00",
         16124 => x"00",
         16125 => x"00",
         16126 => x"00",
         16127 => x"00",
         16128 => x"00",
         16129 => x"00",
         16130 => x"00",
         16131 => x"00",
         16132 => x"00",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"e0",
         18137 => x"cf",
         18138 => x"f9",
         18139 => x"fd",
         18140 => x"c1",
         18141 => x"c5",
         18142 => x"e4",
         18143 => x"ee",
         18144 => x"61",
         18145 => x"65",
         18146 => x"69",
         18147 => x"2a",
         18148 => x"21",
         18149 => x"25",
         18150 => x"29",
         18151 => x"2b",
         18152 => x"01",
         18153 => x"05",
         18154 => x"09",
         18155 => x"0d",
         18156 => x"11",
         18157 => x"15",
         18158 => x"19",
         18159 => x"54",
         18160 => x"81",
         18161 => x"85",
         18162 => x"89",
         18163 => x"8d",
         18164 => x"91",
         18165 => x"95",
         18166 => x"99",
         18167 => x"40",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"02",
         18199 => x"04",
         18200 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"cd",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"e4",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cc",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"ab",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"96",
           269 => x"0b",
           270 => x"0b",
           271 => x"b6",
           272 => x"0b",
           273 => x"0b",
           274 => x"d6",
           275 => x"0b",
           276 => x"0b",
           277 => x"f6",
           278 => x"0b",
           279 => x"0b",
           280 => x"96",
           281 => x"0b",
           282 => x"0b",
           283 => x"b6",
           284 => x"0b",
           285 => x"0b",
           286 => x"d7",
           287 => x"0b",
           288 => x"0b",
           289 => x"f9",
           290 => x"0b",
           291 => x"0b",
           292 => x"9b",
           293 => x"0b",
           294 => x"0b",
           295 => x"bd",
           296 => x"0b",
           297 => x"0b",
           298 => x"df",
           299 => x"0b",
           300 => x"0b",
           301 => x"81",
           302 => x"0b",
           303 => x"0b",
           304 => x"a3",
           305 => x"0b",
           306 => x"0b",
           307 => x"c5",
           308 => x"0b",
           309 => x"0b",
           310 => x"e7",
           311 => x"0b",
           312 => x"0b",
           313 => x"89",
           314 => x"0b",
           315 => x"0b",
           316 => x"ab",
           317 => x"0b",
           318 => x"0b",
           319 => x"cd",
           320 => x"0b",
           321 => x"0b",
           322 => x"ef",
           323 => x"0b",
           324 => x"0b",
           325 => x"91",
           326 => x"0b",
           327 => x"0b",
           328 => x"b3",
           329 => x"0b",
           330 => x"0b",
           331 => x"d5",
           332 => x"0b",
           333 => x"0b",
           334 => x"f7",
           335 => x"0b",
           336 => x"0b",
           337 => x"99",
           338 => x"0b",
           339 => x"0b",
           340 => x"bb",
           341 => x"0b",
           342 => x"0b",
           343 => x"dc",
           344 => x"0b",
           345 => x"0b",
           346 => x"fe",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"90",
           390 => x"f0",
           391 => x"2d",
           392 => x"08",
           393 => x"90",
           394 => x"f0",
           395 => x"2d",
           396 => x"08",
           397 => x"90",
           398 => x"f0",
           399 => x"2d",
           400 => x"08",
           401 => x"90",
           402 => x"f0",
           403 => x"2d",
           404 => x"08",
           405 => x"90",
           406 => x"f0",
           407 => x"2d",
           408 => x"08",
           409 => x"90",
           410 => x"f0",
           411 => x"2d",
           412 => x"08",
           413 => x"90",
           414 => x"f0",
           415 => x"2d",
           416 => x"08",
           417 => x"90",
           418 => x"f0",
           419 => x"2d",
           420 => x"08",
           421 => x"90",
           422 => x"f0",
           423 => x"2d",
           424 => x"08",
           425 => x"90",
           426 => x"f0",
           427 => x"2d",
           428 => x"08",
           429 => x"90",
           430 => x"f0",
           431 => x"2d",
           432 => x"08",
           433 => x"90",
           434 => x"f0",
           435 => x"d1",
           436 => x"f0",
           437 => x"80",
           438 => x"b8",
           439 => x"d5",
           440 => x"b8",
           441 => x"c0",
           442 => x"84",
           443 => x"80",
           444 => x"84",
           445 => x"80",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"90",
           451 => x"f0",
           452 => x"9d",
           453 => x"f0",
           454 => x"80",
           455 => x"b8",
           456 => x"e2",
           457 => x"b8",
           458 => x"c0",
           459 => x"84",
           460 => x"82",
           461 => x"84",
           462 => x"80",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"90",
           468 => x"f0",
           469 => x"8c",
           470 => x"f0",
           471 => x"80",
           472 => x"b8",
           473 => x"fa",
           474 => x"b8",
           475 => x"c0",
           476 => x"84",
           477 => x"82",
           478 => x"84",
           479 => x"80",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"90",
           485 => x"f0",
           486 => x"fa",
           487 => x"f0",
           488 => x"80",
           489 => x"b8",
           490 => x"f3",
           491 => x"b8",
           492 => x"c0",
           493 => x"84",
           494 => x"83",
           495 => x"84",
           496 => x"80",
           497 => x"04",
           498 => x"0c",
           499 => x"2d",
           500 => x"08",
           501 => x"90",
           502 => x"f0",
           503 => x"f5",
           504 => x"f0",
           505 => x"80",
           506 => x"b8",
           507 => x"f5",
           508 => x"b8",
           509 => x"c0",
           510 => x"84",
           511 => x"83",
           512 => x"84",
           513 => x"80",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"90",
           519 => x"f0",
           520 => x"bf",
           521 => x"f0",
           522 => x"80",
           523 => x"b8",
           524 => x"e3",
           525 => x"b8",
           526 => x"c0",
           527 => x"84",
           528 => x"82",
           529 => x"84",
           530 => x"80",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"90",
           536 => x"f0",
           537 => x"89",
           538 => x"f0",
           539 => x"80",
           540 => x"b8",
           541 => x"99",
           542 => x"b8",
           543 => x"c0",
           544 => x"84",
           545 => x"83",
           546 => x"84",
           547 => x"80",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"90",
           553 => x"f0",
           554 => x"81",
           555 => x"f0",
           556 => x"80",
           557 => x"b8",
           558 => x"b9",
           559 => x"b8",
           560 => x"c0",
           561 => x"84",
           562 => x"83",
           563 => x"84",
           564 => x"80",
           565 => x"04",
           566 => x"0c",
           567 => x"2d",
           568 => x"08",
           569 => x"90",
           570 => x"f0",
           571 => x"d1",
           572 => x"f0",
           573 => x"80",
           574 => x"b8",
           575 => x"f5",
           576 => x"b8",
           577 => x"c0",
           578 => x"84",
           579 => x"80",
           580 => x"84",
           581 => x"80",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"90",
           587 => x"f0",
           588 => x"8a",
           589 => x"f0",
           590 => x"80",
           591 => x"b8",
           592 => x"9a",
           593 => x"f0",
           594 => x"80",
           595 => x"b8",
           596 => x"da",
           597 => x"b8",
           598 => x"c0",
           599 => x"84",
           600 => x"81",
           601 => x"84",
           602 => x"80",
           603 => x"04",
           604 => x"0c",
           605 => x"2d",
           606 => x"08",
           607 => x"90",
           608 => x"f0",
           609 => x"80",
           610 => x"f0",
           611 => x"80",
           612 => x"04",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"53",
           621 => x"00",
           622 => x"06",
           623 => x"09",
           624 => x"05",
           625 => x"2b",
           626 => x"06",
           627 => x"04",
           628 => x"72",
           629 => x"05",
           630 => x"05",
           631 => x"72",
           632 => x"53",
           633 => x"51",
           634 => x"04",
           635 => x"70",
           636 => x"27",
           637 => x"71",
           638 => x"53",
           639 => x"0b",
           640 => x"8c",
           641 => x"ce",
           642 => x"fc",
           643 => x"3d",
           644 => x"05",
           645 => x"53",
           646 => x"d4",
           647 => x"81",
           648 => x"3d",
           649 => x"3d",
           650 => x"7c",
           651 => x"81",
           652 => x"80",
           653 => x"56",
           654 => x"80",
           655 => x"2e",
           656 => x"80",
           657 => x"14",
           658 => x"32",
           659 => x"72",
           660 => x"51",
           661 => x"54",
           662 => x"b7",
           663 => x"2e",
           664 => x"51",
           665 => x"84",
           666 => x"53",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"05",
           671 => x"14",
           672 => x"70",
           673 => x"07",
           674 => x"54",
           675 => x"80",
           676 => x"80",
           677 => x"52",
           678 => x"e4",
           679 => x"0d",
           680 => x"84",
           681 => x"88",
           682 => x"f5",
           683 => x"54",
           684 => x"05",
           685 => x"73",
           686 => x"58",
           687 => x"05",
           688 => x"8d",
           689 => x"51",
           690 => x"19",
           691 => x"34",
           692 => x"04",
           693 => x"86",
           694 => x"53",
           695 => x"51",
           696 => x"3d",
           697 => x"3d",
           698 => x"65",
           699 => x"80",
           700 => x"0c",
           701 => x"70",
           702 => x"32",
           703 => x"55",
           704 => x"72",
           705 => x"81",
           706 => x"38",
           707 => x"76",
           708 => x"c5",
           709 => x"7b",
           710 => x"5c",
           711 => x"81",
           712 => x"17",
           713 => x"26",
           714 => x"76",
           715 => x"30",
           716 => x"51",
           717 => x"ae",
           718 => x"2e",
           719 => x"83",
           720 => x"32",
           721 => x"54",
           722 => x"9e",
           723 => x"80",
           724 => x"33",
           725 => x"bd",
           726 => x"08",
           727 => x"b8",
           728 => x"3d",
           729 => x"83",
           730 => x"10",
           731 => x"10",
           732 => x"2b",
           733 => x"19",
           734 => x"0a",
           735 => x"05",
           736 => x"52",
           737 => x"5f",
           738 => x"81",
           739 => x"81",
           740 => x"ff",
           741 => x"7c",
           742 => x"76",
           743 => x"ff",
           744 => x"a5",
           745 => x"06",
           746 => x"73",
           747 => x"5b",
           748 => x"58",
           749 => x"dd",
           750 => x"39",
           751 => x"51",
           752 => x"7b",
           753 => x"fe",
           754 => x"8d",
           755 => x"2a",
           756 => x"54",
           757 => x"38",
           758 => x"06",
           759 => x"95",
           760 => x"53",
           761 => x"26",
           762 => x"10",
           763 => x"f4",
           764 => x"08",
           765 => x"18",
           766 => x"d8",
           767 => x"38",
           768 => x"51",
           769 => x"80",
           770 => x"5b",
           771 => x"38",
           772 => x"80",
           773 => x"f6",
           774 => x"7f",
           775 => x"71",
           776 => x"ff",
           777 => x"58",
           778 => x"b8",
           779 => x"52",
           780 => x"9a",
           781 => x"e4",
           782 => x"06",
           783 => x"08",
           784 => x"56",
           785 => x"26",
           786 => x"b8",
           787 => x"05",
           788 => x"70",
           789 => x"34",
           790 => x"51",
           791 => x"84",
           792 => x"56",
           793 => x"08",
           794 => x"84",
           795 => x"98",
           796 => x"06",
           797 => x"80",
           798 => x"77",
           799 => x"29",
           800 => x"05",
           801 => x"59",
           802 => x"2a",
           803 => x"55",
           804 => x"2e",
           805 => x"84",
           806 => x"f8",
           807 => x"53",
           808 => x"8b",
           809 => x"80",
           810 => x"80",
           811 => x"72",
           812 => x"7a",
           813 => x"81",
           814 => x"72",
           815 => x"38",
           816 => x"70",
           817 => x"54",
           818 => x"24",
           819 => x"7a",
           820 => x"06",
           821 => x"71",
           822 => x"56",
           823 => x"06",
           824 => x"2e",
           825 => x"77",
           826 => x"2b",
           827 => x"7c",
           828 => x"56",
           829 => x"80",
           830 => x"38",
           831 => x"81",
           832 => x"85",
           833 => x"84",
           834 => x"54",
           835 => x"38",
           836 => x"81",
           837 => x"86",
           838 => x"81",
           839 => x"85",
           840 => x"88",
           841 => x"5f",
           842 => x"b2",
           843 => x"84",
           844 => x"fc",
           845 => x"70",
           846 => x"40",
           847 => x"25",
           848 => x"52",
           849 => x"a9",
           850 => x"84",
           851 => x"fc",
           852 => x"70",
           853 => x"40",
           854 => x"24",
           855 => x"81",
           856 => x"80",
           857 => x"78",
           858 => x"0a",
           859 => x"0a",
           860 => x"2c",
           861 => x"80",
           862 => x"38",
           863 => x"51",
           864 => x"78",
           865 => x"0a",
           866 => x"0a",
           867 => x"2c",
           868 => x"74",
           869 => x"38",
           870 => x"70",
           871 => x"55",
           872 => x"81",
           873 => x"80",
           874 => x"d8",
           875 => x"f3",
           876 => x"38",
           877 => x"2e",
           878 => x"7d",
           879 => x"2e",
           880 => x"52",
           881 => x"33",
           882 => x"a5",
           883 => x"b8",
           884 => x"81",
           885 => x"74",
           886 => x"7a",
           887 => x"a7",
           888 => x"84",
           889 => x"fc",
           890 => x"70",
           891 => x"40",
           892 => x"25",
           893 => x"7c",
           894 => x"86",
           895 => x"39",
           896 => x"5b",
           897 => x"7c",
           898 => x"76",
           899 => x"fa",
           900 => x"80",
           901 => x"80",
           902 => x"60",
           903 => x"71",
           904 => x"ff",
           905 => x"59",
           906 => x"fb",
           907 => x"60",
           908 => x"fe",
           909 => x"83",
           910 => x"98",
           911 => x"7c",
           912 => x"29",
           913 => x"05",
           914 => x"5e",
           915 => x"57",
           916 => x"87",
           917 => x"06",
           918 => x"fe",
           919 => x"78",
           920 => x"29",
           921 => x"05",
           922 => x"5a",
           923 => x"7f",
           924 => x"38",
           925 => x"51",
           926 => x"e2",
           927 => x"70",
           928 => x"06",
           929 => x"83",
           930 => x"fe",
           931 => x"52",
           932 => x"05",
           933 => x"85",
           934 => x"39",
           935 => x"83",
           936 => x"5b",
           937 => x"ff",
           938 => x"ab",
           939 => x"75",
           940 => x"57",
           941 => x"b9",
           942 => x"75",
           943 => x"81",
           944 => x"78",
           945 => x"29",
           946 => x"05",
           947 => x"5a",
           948 => x"e3",
           949 => x"70",
           950 => x"56",
           951 => x"c6",
           952 => x"39",
           953 => x"05",
           954 => x"53",
           955 => x"80",
           956 => x"df",
           957 => x"ff",
           958 => x"84",
           959 => x"fa",
           960 => x"84",
           961 => x"58",
           962 => x"89",
           963 => x"39",
           964 => x"5b",
           965 => x"58",
           966 => x"f9",
           967 => x"39",
           968 => x"05",
           969 => x"81",
           970 => x"41",
           971 => x"8a",
           972 => x"87",
           973 => x"b8",
           974 => x"ff",
           975 => x"71",
           976 => x"54",
           977 => x"2c",
           978 => x"39",
           979 => x"07",
           980 => x"5b",
           981 => x"38",
           982 => x"7f",
           983 => x"71",
           984 => x"06",
           985 => x"54",
           986 => x"38",
           987 => x"bb",
           988 => x"e4",
           989 => x"ff",
           990 => x"31",
           991 => x"5a",
           992 => x"81",
           993 => x"33",
           994 => x"f7",
           995 => x"c9",
           996 => x"84",
           997 => x"fc",
           998 => x"70",
           999 => x"54",
          1000 => x"25",
          1001 => x"7c",
          1002 => x"83",
          1003 => x"39",
          1004 => x"51",
          1005 => x"79",
          1006 => x"81",
          1007 => x"38",
          1008 => x"51",
          1009 => x"7a",
          1010 => x"06",
          1011 => x"2e",
          1012 => x"fa",
          1013 => x"98",
          1014 => x"31",
          1015 => x"90",
          1016 => x"80",
          1017 => x"51",
          1018 => x"90",
          1019 => x"39",
          1020 => x"51",
          1021 => x"7e",
          1022 => x"73",
          1023 => x"a2",
          1024 => x"39",
          1025 => x"98",
          1026 => x"e5",
          1027 => x"06",
          1028 => x"2e",
          1029 => x"fb",
          1030 => x"74",
          1031 => x"70",
          1032 => x"53",
          1033 => x"7c",
          1034 => x"82",
          1035 => x"39",
          1036 => x"51",
          1037 => x"ff",
          1038 => x"52",
          1039 => x"8b",
          1040 => x"e4",
          1041 => x"ff",
          1042 => x"31",
          1043 => x"5a",
          1044 => x"7a",
          1045 => x"30",
          1046 => x"bf",
          1047 => x"5b",
          1048 => x"fe",
          1049 => x"d4",
          1050 => x"75",
          1051 => x"f3",
          1052 => x"3d",
          1053 => x"3d",
          1054 => x"80",
          1055 => x"c8",
          1056 => x"33",
          1057 => x"81",
          1058 => x"06",
          1059 => x"55",
          1060 => x"72",
          1061 => x"81",
          1062 => x"38",
          1063 => x"05",
          1064 => x"72",
          1065 => x"38",
          1066 => x"08",
          1067 => x"90",
          1068 => x"72",
          1069 => x"e4",
          1070 => x"83",
          1071 => x"74",
          1072 => x"56",
          1073 => x"80",
          1074 => x"84",
          1075 => x"54",
          1076 => x"d4",
          1077 => x"84",
          1078 => x"52",
          1079 => x"14",
          1080 => x"2d",
          1081 => x"08",
          1082 => x"38",
          1083 => x"56",
          1084 => x"e4",
          1085 => x"0d",
          1086 => x"0d",
          1087 => x"54",
          1088 => x"16",
          1089 => x"2a",
          1090 => x"81",
          1091 => x"57",
          1092 => x"72",
          1093 => x"81",
          1094 => x"73",
          1095 => x"55",
          1096 => x"77",
          1097 => x"06",
          1098 => x"56",
          1099 => x"e4",
          1100 => x"0d",
          1101 => x"81",
          1102 => x"53",
          1103 => x"ea",
          1104 => x"72",
          1105 => x"08",
          1106 => x"84",
          1107 => x"80",
          1108 => x"ff",
          1109 => x"05",
          1110 => x"57",
          1111 => x"ca",
          1112 => x"0d",
          1113 => x"08",
          1114 => x"85",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"11",
          1118 => x"2a",
          1119 => x"06",
          1120 => x"57",
          1121 => x"ae",
          1122 => x"2a",
          1123 => x"73",
          1124 => x"38",
          1125 => x"53",
          1126 => x"08",
          1127 => x"74",
          1128 => x"76",
          1129 => x"81",
          1130 => x"8c",
          1131 => x"81",
          1132 => x"0c",
          1133 => x"84",
          1134 => x"88",
          1135 => x"74",
          1136 => x"ff",
          1137 => x"15",
          1138 => x"2d",
          1139 => x"b8",
          1140 => x"38",
          1141 => x"81",
          1142 => x"0c",
          1143 => x"39",
          1144 => x"77",
          1145 => x"70",
          1146 => x"70",
          1147 => x"06",
          1148 => x"56",
          1149 => x"b3",
          1150 => x"2a",
          1151 => x"71",
          1152 => x"82",
          1153 => x"52",
          1154 => x"80",
          1155 => x"08",
          1156 => x"53",
          1157 => x"80",
          1158 => x"13",
          1159 => x"16",
          1160 => x"8c",
          1161 => x"81",
          1162 => x"73",
          1163 => x"0c",
          1164 => x"04",
          1165 => x"06",
          1166 => x"17",
          1167 => x"08",
          1168 => x"17",
          1169 => x"33",
          1170 => x"0c",
          1171 => x"04",
          1172 => x"16",
          1173 => x"2d",
          1174 => x"08",
          1175 => x"e4",
          1176 => x"ff",
          1177 => x"16",
          1178 => x"07",
          1179 => x"b8",
          1180 => x"2e",
          1181 => x"a0",
          1182 => x"85",
          1183 => x"54",
          1184 => x"e4",
          1185 => x"0d",
          1186 => x"07",
          1187 => x"17",
          1188 => x"ec",
          1189 => x"0d",
          1190 => x"54",
          1191 => x"70",
          1192 => x"33",
          1193 => x"38",
          1194 => x"72",
          1195 => x"54",
          1196 => x"72",
          1197 => x"54",
          1198 => x"38",
          1199 => x"e4",
          1200 => x"0d",
          1201 => x"0d",
          1202 => x"7a",
          1203 => x"54",
          1204 => x"9d",
          1205 => x"27",
          1206 => x"80",
          1207 => x"71",
          1208 => x"53",
          1209 => x"81",
          1210 => x"ff",
          1211 => x"ef",
          1212 => x"b8",
          1213 => x"3d",
          1214 => x"12",
          1215 => x"27",
          1216 => x"14",
          1217 => x"ff",
          1218 => x"53",
          1219 => x"73",
          1220 => x"51",
          1221 => x"d9",
          1222 => x"ff",
          1223 => x"71",
          1224 => x"ff",
          1225 => x"df",
          1226 => x"fe",
          1227 => x"70",
          1228 => x"70",
          1229 => x"33",
          1230 => x"38",
          1231 => x"74",
          1232 => x"e4",
          1233 => x"3d",
          1234 => x"3d",
          1235 => x"71",
          1236 => x"72",
          1237 => x"54",
          1238 => x"72",
          1239 => x"54",
          1240 => x"38",
          1241 => x"e4",
          1242 => x"0d",
          1243 => x"0d",
          1244 => x"79",
          1245 => x"54",
          1246 => x"93",
          1247 => x"81",
          1248 => x"73",
          1249 => x"55",
          1250 => x"51",
          1251 => x"73",
          1252 => x"0c",
          1253 => x"04",
          1254 => x"76",
          1255 => x"56",
          1256 => x"2e",
          1257 => x"33",
          1258 => x"05",
          1259 => x"52",
          1260 => x"09",
          1261 => x"38",
          1262 => x"71",
          1263 => x"38",
          1264 => x"72",
          1265 => x"51",
          1266 => x"e4",
          1267 => x"0d",
          1268 => x"2e",
          1269 => x"33",
          1270 => x"72",
          1271 => x"38",
          1272 => x"52",
          1273 => x"80",
          1274 => x"72",
          1275 => x"b8",
          1276 => x"3d",
          1277 => x"84",
          1278 => x"86",
          1279 => x"fb",
          1280 => x"79",
          1281 => x"56",
          1282 => x"84",
          1283 => x"84",
          1284 => x"81",
          1285 => x"81",
          1286 => x"84",
          1287 => x"54",
          1288 => x"08",
          1289 => x"38",
          1290 => x"08",
          1291 => x"74",
          1292 => x"75",
          1293 => x"e4",
          1294 => x"b1",
          1295 => x"e4",
          1296 => x"84",
          1297 => x"87",
          1298 => x"fd",
          1299 => x"77",
          1300 => x"55",
          1301 => x"80",
          1302 => x"72",
          1303 => x"54",
          1304 => x"80",
          1305 => x"ff",
          1306 => x"ff",
          1307 => x"06",
          1308 => x"13",
          1309 => x"52",
          1310 => x"b8",
          1311 => x"3d",
          1312 => x"3d",
          1313 => x"79",
          1314 => x"54",
          1315 => x"2e",
          1316 => x"72",
          1317 => x"54",
          1318 => x"51",
          1319 => x"73",
          1320 => x"0c",
          1321 => x"04",
          1322 => x"78",
          1323 => x"a0",
          1324 => x"2e",
          1325 => x"51",
          1326 => x"84",
          1327 => x"52",
          1328 => x"73",
          1329 => x"38",
          1330 => x"e3",
          1331 => x"b8",
          1332 => x"53",
          1333 => x"9f",
          1334 => x"38",
          1335 => x"9f",
          1336 => x"38",
          1337 => x"71",
          1338 => x"31",
          1339 => x"57",
          1340 => x"80",
          1341 => x"2e",
          1342 => x"10",
          1343 => x"07",
          1344 => x"07",
          1345 => x"ff",
          1346 => x"70",
          1347 => x"72",
          1348 => x"31",
          1349 => x"56",
          1350 => x"58",
          1351 => x"da",
          1352 => x"76",
          1353 => x"84",
          1354 => x"88",
          1355 => x"fc",
          1356 => x"70",
          1357 => x"06",
          1358 => x"72",
          1359 => x"70",
          1360 => x"71",
          1361 => x"2a",
          1362 => x"80",
          1363 => x"70",
          1364 => x"2b",
          1365 => x"74",
          1366 => x"81",
          1367 => x"30",
          1368 => x"82",
          1369 => x"31",
          1370 => x"55",
          1371 => x"05",
          1372 => x"70",
          1373 => x"25",
          1374 => x"31",
          1375 => x"70",
          1376 => x"32",
          1377 => x"70",
          1378 => x"31",
          1379 => x"05",
          1380 => x"0c",
          1381 => x"55",
          1382 => x"5a",
          1383 => x"55",
          1384 => x"56",
          1385 => x"56",
          1386 => x"3d",
          1387 => x"3d",
          1388 => x"70",
          1389 => x"54",
          1390 => x"3f",
          1391 => x"08",
          1392 => x"71",
          1393 => x"e4",
          1394 => x"3d",
          1395 => x"3d",
          1396 => x"58",
          1397 => x"76",
          1398 => x"38",
          1399 => x"cf",
          1400 => x"e4",
          1401 => x"13",
          1402 => x"2e",
          1403 => x"51",
          1404 => x"72",
          1405 => x"08",
          1406 => x"53",
          1407 => x"80",
          1408 => x"53",
          1409 => x"be",
          1410 => x"74",
          1411 => x"72",
          1412 => x"2b",
          1413 => x"55",
          1414 => x"76",
          1415 => x"72",
          1416 => x"2a",
          1417 => x"77",
          1418 => x"31",
          1419 => x"2c",
          1420 => x"7b",
          1421 => x"71",
          1422 => x"5c",
          1423 => x"55",
          1424 => x"74",
          1425 => x"84",
          1426 => x"88",
          1427 => x"fa",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"7b",
          1431 => x"2c",
          1432 => x"73",
          1433 => x"31",
          1434 => x"31",
          1435 => x"59",
          1436 => x"b4",
          1437 => x"e4",
          1438 => x"75",
          1439 => x"e4",
          1440 => x"0d",
          1441 => x"0d",
          1442 => x"57",
          1443 => x"0c",
          1444 => x"33",
          1445 => x"73",
          1446 => x"81",
          1447 => x"81",
          1448 => x"0c",
          1449 => x"55",
          1450 => x"f3",
          1451 => x"2e",
          1452 => x"73",
          1453 => x"83",
          1454 => x"58",
          1455 => x"89",
          1456 => x"38",
          1457 => x"56",
          1458 => x"80",
          1459 => x"e0",
          1460 => x"38",
          1461 => x"81",
          1462 => x"53",
          1463 => x"81",
          1464 => x"53",
          1465 => x"8f",
          1466 => x"70",
          1467 => x"54",
          1468 => x"27",
          1469 => x"72",
          1470 => x"83",
          1471 => x"29",
          1472 => x"70",
          1473 => x"33",
          1474 => x"73",
          1475 => x"be",
          1476 => x"2e",
          1477 => x"30",
          1478 => x"0c",
          1479 => x"84",
          1480 => x"8b",
          1481 => x"81",
          1482 => x"79",
          1483 => x"56",
          1484 => x"b0",
          1485 => x"06",
          1486 => x"81",
          1487 => x"0c",
          1488 => x"55",
          1489 => x"2e",
          1490 => x"58",
          1491 => x"2e",
          1492 => x"56",
          1493 => x"c6",
          1494 => x"53",
          1495 => x"58",
          1496 => x"fe",
          1497 => x"84",
          1498 => x"8b",
          1499 => x"82",
          1500 => x"70",
          1501 => x"33",
          1502 => x"56",
          1503 => x"80",
          1504 => x"e4",
          1505 => x"0d",
          1506 => x"0d",
          1507 => x"57",
          1508 => x"0c",
          1509 => x"33",
          1510 => x"73",
          1511 => x"81",
          1512 => x"81",
          1513 => x"0c",
          1514 => x"55",
          1515 => x"f3",
          1516 => x"2e",
          1517 => x"73",
          1518 => x"83",
          1519 => x"58",
          1520 => x"89",
          1521 => x"38",
          1522 => x"56",
          1523 => x"80",
          1524 => x"e0",
          1525 => x"38",
          1526 => x"81",
          1527 => x"53",
          1528 => x"81",
          1529 => x"53",
          1530 => x"8f",
          1531 => x"70",
          1532 => x"54",
          1533 => x"27",
          1534 => x"72",
          1535 => x"83",
          1536 => x"29",
          1537 => x"70",
          1538 => x"33",
          1539 => x"73",
          1540 => x"be",
          1541 => x"2e",
          1542 => x"30",
          1543 => x"0c",
          1544 => x"84",
          1545 => x"8b",
          1546 => x"81",
          1547 => x"79",
          1548 => x"56",
          1549 => x"b0",
          1550 => x"06",
          1551 => x"81",
          1552 => x"0c",
          1553 => x"55",
          1554 => x"2e",
          1555 => x"58",
          1556 => x"2e",
          1557 => x"56",
          1558 => x"c6",
          1559 => x"53",
          1560 => x"58",
          1561 => x"fe",
          1562 => x"84",
          1563 => x"8b",
          1564 => x"82",
          1565 => x"70",
          1566 => x"33",
          1567 => x"56",
          1568 => x"80",
          1569 => x"e4",
          1570 => x"0d",
          1571 => x"d1",
          1572 => x"e4",
          1573 => x"06",
          1574 => x"0c",
          1575 => x"0d",
          1576 => x"93",
          1577 => x"71",
          1578 => x"bd",
          1579 => x"71",
          1580 => x"ce",
          1581 => x"be",
          1582 => x"0d",
          1583 => x"9c",
          1584 => x"3f",
          1585 => x"04",
          1586 => x"51",
          1587 => x"83",
          1588 => x"83",
          1589 => x"ef",
          1590 => x"3d",
          1591 => x"ce",
          1592 => x"92",
          1593 => x"0d",
          1594 => x"f4",
          1595 => x"3f",
          1596 => x"04",
          1597 => x"51",
          1598 => x"83",
          1599 => x"83",
          1600 => x"ee",
          1601 => x"3d",
          1602 => x"cf",
          1603 => x"e6",
          1604 => x"0d",
          1605 => x"e0",
          1606 => x"3f",
          1607 => x"04",
          1608 => x"51",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ee",
          1612 => x"3d",
          1613 => x"d0",
          1614 => x"ba",
          1615 => x"0d",
          1616 => x"c4",
          1617 => x"3f",
          1618 => x"04",
          1619 => x"51",
          1620 => x"83",
          1621 => x"83",
          1622 => x"ee",
          1623 => x"3d",
          1624 => x"d0",
          1625 => x"8e",
          1626 => x"0d",
          1627 => x"88",
          1628 => x"3f",
          1629 => x"04",
          1630 => x"51",
          1631 => x"83",
          1632 => x"83",
          1633 => x"ed",
          1634 => x"3d",
          1635 => x"d1",
          1636 => x"e2",
          1637 => x"0d",
          1638 => x"0d",
          1639 => x"05",
          1640 => x"33",
          1641 => x"68",
          1642 => x"7b",
          1643 => x"51",
          1644 => x"78",
          1645 => x"ff",
          1646 => x"81",
          1647 => x"07",
          1648 => x"06",
          1649 => x"57",
          1650 => x"38",
          1651 => x"52",
          1652 => x"52",
          1653 => x"c8",
          1654 => x"e4",
          1655 => x"b8",
          1656 => x"2e",
          1657 => x"77",
          1658 => x"86",
          1659 => x"70",
          1660 => x"25",
          1661 => x"9f",
          1662 => x"53",
          1663 => x"77",
          1664 => x"38",
          1665 => x"88",
          1666 => x"87",
          1667 => x"e0",
          1668 => x"78",
          1669 => x"51",
          1670 => x"84",
          1671 => x"54",
          1672 => x"53",
          1673 => x"d1",
          1674 => x"df",
          1675 => x"b8",
          1676 => x"3d",
          1677 => x"b8",
          1678 => x"c0",
          1679 => x"84",
          1680 => x"59",
          1681 => x"05",
          1682 => x"53",
          1683 => x"51",
          1684 => x"3f",
          1685 => x"08",
          1686 => x"e4",
          1687 => x"38",
          1688 => x"80",
          1689 => x"38",
          1690 => x"17",
          1691 => x"39",
          1692 => x"74",
          1693 => x"3f",
          1694 => x"08",
          1695 => x"f4",
          1696 => x"b8",
          1697 => x"83",
          1698 => x"78",
          1699 => x"c0",
          1700 => x"3f",
          1701 => x"f8",
          1702 => x"02",
          1703 => x"05",
          1704 => x"ff",
          1705 => x"7b",
          1706 => x"fd",
          1707 => x"b8",
          1708 => x"38",
          1709 => x"91",
          1710 => x"2e",
          1711 => x"84",
          1712 => x"8a",
          1713 => x"78",
          1714 => x"c4",
          1715 => x"60",
          1716 => x"e4",
          1717 => x"7e",
          1718 => x"84",
          1719 => x"84",
          1720 => x"8a",
          1721 => x"f3",
          1722 => x"61",
          1723 => x"05",
          1724 => x"33",
          1725 => x"68",
          1726 => x"5c",
          1727 => x"78",
          1728 => x"82",
          1729 => x"83",
          1730 => x"dd",
          1731 => x"d1",
          1732 => x"f7",
          1733 => x"73",
          1734 => x"38",
          1735 => x"81",
          1736 => x"a0",
          1737 => x"38",
          1738 => x"72",
          1739 => x"a7",
          1740 => x"52",
          1741 => x"51",
          1742 => x"81",
          1743 => x"c8",
          1744 => x"a0",
          1745 => x"3f",
          1746 => x"dc",
          1747 => x"80",
          1748 => x"3f",
          1749 => x"79",
          1750 => x"38",
          1751 => x"33",
          1752 => x"55",
          1753 => x"83",
          1754 => x"80",
          1755 => x"27",
          1756 => x"53",
          1757 => x"70",
          1758 => x"56",
          1759 => x"2e",
          1760 => x"fe",
          1761 => x"ee",
          1762 => x"c8",
          1763 => x"51",
          1764 => x"81",
          1765 => x"76",
          1766 => x"83",
          1767 => x"e9",
          1768 => x"18",
          1769 => x"58",
          1770 => x"a8",
          1771 => x"e4",
          1772 => x"70",
          1773 => x"54",
          1774 => x"81",
          1775 => x"9b",
          1776 => x"38",
          1777 => x"76",
          1778 => x"b9",
          1779 => x"84",
          1780 => x"8f",
          1781 => x"83",
          1782 => x"dc",
          1783 => x"14",
          1784 => x"08",
          1785 => x"51",
          1786 => x"78",
          1787 => x"b8",
          1788 => x"39",
          1789 => x"51",
          1790 => x"82",
          1791 => x"c8",
          1792 => x"a0",
          1793 => x"3f",
          1794 => x"fe",
          1795 => x"18",
          1796 => x"27",
          1797 => x"22",
          1798 => x"8c",
          1799 => x"3f",
          1800 => x"d4",
          1801 => x"54",
          1802 => x"c5",
          1803 => x"26",
          1804 => x"99",
          1805 => x"94",
          1806 => x"3f",
          1807 => x"d4",
          1808 => x"54",
          1809 => x"a9",
          1810 => x"27",
          1811 => x"73",
          1812 => x"7a",
          1813 => x"72",
          1814 => x"d1",
          1815 => x"ab",
          1816 => x"84",
          1817 => x"53",
          1818 => x"ea",
          1819 => x"74",
          1820 => x"fd",
          1821 => x"d4",
          1822 => x"73",
          1823 => x"3f",
          1824 => x"fe",
          1825 => x"ce",
          1826 => x"b8",
          1827 => x"ff",
          1828 => x"59",
          1829 => x"fc",
          1830 => x"59",
          1831 => x"2e",
          1832 => x"fc",
          1833 => x"59",
          1834 => x"80",
          1835 => x"3f",
          1836 => x"08",
          1837 => x"98",
          1838 => x"32",
          1839 => x"9b",
          1840 => x"70",
          1841 => x"75",
          1842 => x"55",
          1843 => x"58",
          1844 => x"25",
          1845 => x"80",
          1846 => x"3f",
          1847 => x"08",
          1848 => x"98",
          1849 => x"32",
          1850 => x"9b",
          1851 => x"70",
          1852 => x"75",
          1853 => x"55",
          1854 => x"58",
          1855 => x"24",
          1856 => x"fd",
          1857 => x"0b",
          1858 => x"0c",
          1859 => x"04",
          1860 => x"87",
          1861 => x"08",
          1862 => x"3f",
          1863 => x"ed",
          1864 => x"dc",
          1865 => x"3f",
          1866 => x"e1",
          1867 => x"2a",
          1868 => x"51",
          1869 => x"b7",
          1870 => x"2a",
          1871 => x"51",
          1872 => x"89",
          1873 => x"2a",
          1874 => x"51",
          1875 => x"db",
          1876 => x"2a",
          1877 => x"51",
          1878 => x"ad",
          1879 => x"2a",
          1880 => x"51",
          1881 => x"ff",
          1882 => x"2a",
          1883 => x"51",
          1884 => x"d2",
          1885 => x"2a",
          1886 => x"51",
          1887 => x"38",
          1888 => x"81",
          1889 => x"88",
          1890 => x"3f",
          1891 => x"04",
          1892 => x"f9",
          1893 => x"f4",
          1894 => x"3f",
          1895 => x"ed",
          1896 => x"3f",
          1897 => x"04",
          1898 => x"e1",
          1899 => x"88",
          1900 => x"3f",
          1901 => x"d5",
          1902 => x"2a",
          1903 => x"72",
          1904 => x"38",
          1905 => x"51",
          1906 => x"83",
          1907 => x"9b",
          1908 => x"51",
          1909 => x"72",
          1910 => x"81",
          1911 => x"71",
          1912 => x"9c",
          1913 => x"81",
          1914 => x"3f",
          1915 => x"51",
          1916 => x"80",
          1917 => x"3f",
          1918 => x"70",
          1919 => x"52",
          1920 => x"fe",
          1921 => x"be",
          1922 => x"9b",
          1923 => x"d3",
          1924 => x"91",
          1925 => x"9a",
          1926 => x"85",
          1927 => x"06",
          1928 => x"80",
          1929 => x"38",
          1930 => x"81",
          1931 => x"3f",
          1932 => x"51",
          1933 => x"80",
          1934 => x"3f",
          1935 => x"70",
          1936 => x"52",
          1937 => x"fe",
          1938 => x"bd",
          1939 => x"9a",
          1940 => x"d3",
          1941 => x"cd",
          1942 => x"9a",
          1943 => x"83",
          1944 => x"06",
          1945 => x"80",
          1946 => x"38",
          1947 => x"81",
          1948 => x"3f",
          1949 => x"51",
          1950 => x"80",
          1951 => x"3f",
          1952 => x"70",
          1953 => x"52",
          1954 => x"fd",
          1955 => x"bd",
          1956 => x"0d",
          1957 => x"41",
          1958 => x"cf",
          1959 => x"81",
          1960 => x"81",
          1961 => x"84",
          1962 => x"81",
          1963 => x"3d",
          1964 => x"61",
          1965 => x"38",
          1966 => x"51",
          1967 => x"98",
          1968 => x"d5",
          1969 => x"c3",
          1970 => x"80",
          1971 => x"52",
          1972 => x"ae",
          1973 => x"83",
          1974 => x"70",
          1975 => x"5b",
          1976 => x"2e",
          1977 => x"79",
          1978 => x"88",
          1979 => x"ff",
          1980 => x"82",
          1981 => x"38",
          1982 => x"5a",
          1983 => x"83",
          1984 => x"33",
          1985 => x"2e",
          1986 => x"8c",
          1987 => x"70",
          1988 => x"7b",
          1989 => x"38",
          1990 => x"9b",
          1991 => x"7b",
          1992 => x"ed",
          1993 => x"08",
          1994 => x"ff",
          1995 => x"e4",
          1996 => x"e4",
          1997 => x"53",
          1998 => x"5d",
          1999 => x"84",
          2000 => x"8b",
          2001 => x"33",
          2002 => x"2e",
          2003 => x"81",
          2004 => x"ff",
          2005 => x"9b",
          2006 => x"38",
          2007 => x"5c",
          2008 => x"fe",
          2009 => x"f8",
          2010 => x"e9",
          2011 => x"b8",
          2012 => x"84",
          2013 => x"80",
          2014 => x"38",
          2015 => x"08",
          2016 => x"ff",
          2017 => x"91",
          2018 => x"b8",
          2019 => x"62",
          2020 => x"7a",
          2021 => x"84",
          2022 => x"e4",
          2023 => x"8b",
          2024 => x"e4",
          2025 => x"80",
          2026 => x"0b",
          2027 => x"5b",
          2028 => x"8d",
          2029 => x"82",
          2030 => x"38",
          2031 => x"82",
          2032 => x"54",
          2033 => x"d5",
          2034 => x"51",
          2035 => x"83",
          2036 => x"84",
          2037 => x"7d",
          2038 => x"80",
          2039 => x"0a",
          2040 => x"0a",
          2041 => x"f5",
          2042 => x"b8",
          2043 => x"b8",
          2044 => x"70",
          2045 => x"07",
          2046 => x"5b",
          2047 => x"5a",
          2048 => x"83",
          2049 => x"78",
          2050 => x"78",
          2051 => x"38",
          2052 => x"81",
          2053 => x"5a",
          2054 => x"38",
          2055 => x"61",
          2056 => x"5d",
          2057 => x"38",
          2058 => x"81",
          2059 => x"51",
          2060 => x"3f",
          2061 => x"51",
          2062 => x"7e",
          2063 => x"53",
          2064 => x"51",
          2065 => x"0b",
          2066 => x"d8",
          2067 => x"ff",
          2068 => x"79",
          2069 => x"81",
          2070 => x"b4",
          2071 => x"f4",
          2072 => x"bc",
          2073 => x"e4",
          2074 => x"38",
          2075 => x"0b",
          2076 => x"34",
          2077 => x"53",
          2078 => x"7e",
          2079 => x"b7",
          2080 => x"e4",
          2081 => x"a0",
          2082 => x"e4",
          2083 => x"e6",
          2084 => x"83",
          2085 => x"70",
          2086 => x"5f",
          2087 => x"2e",
          2088 => x"fc",
          2089 => x"39",
          2090 => x"51",
          2091 => x"3f",
          2092 => x"0b",
          2093 => x"34",
          2094 => x"53",
          2095 => x"7e",
          2096 => x"3f",
          2097 => x"5a",
          2098 => x"38",
          2099 => x"1a",
          2100 => x"1b",
          2101 => x"81",
          2102 => x"80",
          2103 => x"10",
          2104 => x"05",
          2105 => x"04",
          2106 => x"d5",
          2107 => x"51",
          2108 => x"60",
          2109 => x"84",
          2110 => x"82",
          2111 => x"84",
          2112 => x"61",
          2113 => x"06",
          2114 => x"81",
          2115 => x"45",
          2116 => x"ae",
          2117 => x"98",
          2118 => x"3f",
          2119 => x"92",
          2120 => x"90",
          2121 => x"a8",
          2122 => x"83",
          2123 => x"80",
          2124 => x"b0",
          2125 => x"d2",
          2126 => x"93",
          2127 => x"9a",
          2128 => x"39",
          2129 => x"fa",
          2130 => x"52",
          2131 => x"93",
          2132 => x"39",
          2133 => x"3f",
          2134 => x"83",
          2135 => x"de",
          2136 => x"59",
          2137 => x"d5",
          2138 => x"8a",
          2139 => x"3f",
          2140 => x"b8",
          2141 => x"11",
          2142 => x"05",
          2143 => x"3f",
          2144 => x"08",
          2145 => x"ba",
          2146 => x"83",
          2147 => x"d0",
          2148 => x"5a",
          2149 => x"b8",
          2150 => x"2e",
          2151 => x"84",
          2152 => x"52",
          2153 => x"51",
          2154 => x"fa",
          2155 => x"3d",
          2156 => x"53",
          2157 => x"51",
          2158 => x"84",
          2159 => x"80",
          2160 => x"38",
          2161 => x"d6",
          2162 => x"bf",
          2163 => x"78",
          2164 => x"fe",
          2165 => x"ff",
          2166 => x"e9",
          2167 => x"b8",
          2168 => x"2e",
          2169 => x"b8",
          2170 => x"11",
          2171 => x"05",
          2172 => x"3f",
          2173 => x"08",
          2174 => x"64",
          2175 => x"53",
          2176 => x"d6",
          2177 => x"83",
          2178 => x"c4",
          2179 => x"f8",
          2180 => x"d0",
          2181 => x"48",
          2182 => x"78",
          2183 => x"a2",
          2184 => x"26",
          2185 => x"64",
          2186 => x"46",
          2187 => x"b8",
          2188 => x"11",
          2189 => x"05",
          2190 => x"3f",
          2191 => x"08",
          2192 => x"fe",
          2193 => x"fe",
          2194 => x"ff",
          2195 => x"e8",
          2196 => x"b8",
          2197 => x"b0",
          2198 => x"78",
          2199 => x"52",
          2200 => x"51",
          2201 => x"84",
          2202 => x"53",
          2203 => x"7e",
          2204 => x"3f",
          2205 => x"33",
          2206 => x"2e",
          2207 => x"78",
          2208 => x"ca",
          2209 => x"05",
          2210 => x"cf",
          2211 => x"ff",
          2212 => x"ff",
          2213 => x"e9",
          2214 => x"b8",
          2215 => x"2e",
          2216 => x"b8",
          2217 => x"11",
          2218 => x"05",
          2219 => x"3f",
          2220 => x"08",
          2221 => x"8a",
          2222 => x"fe",
          2223 => x"ff",
          2224 => x"e9",
          2225 => x"b8",
          2226 => x"2e",
          2227 => x"83",
          2228 => x"ce",
          2229 => x"67",
          2230 => x"7c",
          2231 => x"38",
          2232 => x"7a",
          2233 => x"5a",
          2234 => x"95",
          2235 => x"79",
          2236 => x"53",
          2237 => x"d6",
          2238 => x"8f",
          2239 => x"5b",
          2240 => x"81",
          2241 => x"d2",
          2242 => x"ff",
          2243 => x"ff",
          2244 => x"e8",
          2245 => x"b8",
          2246 => x"2e",
          2247 => x"b8",
          2248 => x"11",
          2249 => x"05",
          2250 => x"3f",
          2251 => x"08",
          2252 => x"8e",
          2253 => x"fe",
          2254 => x"ff",
          2255 => x"e8",
          2256 => x"b8",
          2257 => x"2e",
          2258 => x"83",
          2259 => x"cd",
          2260 => x"5a",
          2261 => x"82",
          2262 => x"5c",
          2263 => x"05",
          2264 => x"34",
          2265 => x"46",
          2266 => x"3d",
          2267 => x"53",
          2268 => x"51",
          2269 => x"84",
          2270 => x"80",
          2271 => x"38",
          2272 => x"fc",
          2273 => x"80",
          2274 => x"fd",
          2275 => x"e4",
          2276 => x"68",
          2277 => x"52",
          2278 => x"51",
          2279 => x"84",
          2280 => x"53",
          2281 => x"7e",
          2282 => x"3f",
          2283 => x"33",
          2284 => x"2e",
          2285 => x"78",
          2286 => x"97",
          2287 => x"05",
          2288 => x"68",
          2289 => x"db",
          2290 => x"34",
          2291 => x"49",
          2292 => x"fc",
          2293 => x"80",
          2294 => x"ad",
          2295 => x"e4",
          2296 => x"f5",
          2297 => x"59",
          2298 => x"05",
          2299 => x"68",
          2300 => x"b8",
          2301 => x"11",
          2302 => x"05",
          2303 => x"3f",
          2304 => x"08",
          2305 => x"f5",
          2306 => x"3d",
          2307 => x"53",
          2308 => x"51",
          2309 => x"84",
          2310 => x"80",
          2311 => x"38",
          2312 => x"fc",
          2313 => x"80",
          2314 => x"dd",
          2315 => x"e4",
          2316 => x"f5",
          2317 => x"3d",
          2318 => x"53",
          2319 => x"51",
          2320 => x"84",
          2321 => x"86",
          2322 => x"e4",
          2323 => x"d7",
          2324 => x"b7",
          2325 => x"5b",
          2326 => x"27",
          2327 => x"5b",
          2328 => x"84",
          2329 => x"79",
          2330 => x"38",
          2331 => x"f1",
          2332 => x"39",
          2333 => x"80",
          2334 => x"96",
          2335 => x"e4",
          2336 => x"ff",
          2337 => x"59",
          2338 => x"81",
          2339 => x"e4",
          2340 => x"51",
          2341 => x"84",
          2342 => x"80",
          2343 => x"38",
          2344 => x"08",
          2345 => x"3f",
          2346 => x"b8",
          2347 => x"11",
          2348 => x"05",
          2349 => x"3f",
          2350 => x"08",
          2351 => x"f1",
          2352 => x"79",
          2353 => x"c0",
          2354 => x"a0",
          2355 => x"3d",
          2356 => x"53",
          2357 => x"51",
          2358 => x"84",
          2359 => x"91",
          2360 => x"e8",
          2361 => x"80",
          2362 => x"38",
          2363 => x"08",
          2364 => x"fe",
          2365 => x"ff",
          2366 => x"e5",
          2367 => x"b8",
          2368 => x"2e",
          2369 => x"66",
          2370 => x"88",
          2371 => x"81",
          2372 => x"32",
          2373 => x"72",
          2374 => x"7e",
          2375 => x"5d",
          2376 => x"88",
          2377 => x"2e",
          2378 => x"46",
          2379 => x"51",
          2380 => x"80",
          2381 => x"65",
          2382 => x"68",
          2383 => x"3f",
          2384 => x"51",
          2385 => x"f2",
          2386 => x"64",
          2387 => x"64",
          2388 => x"b8",
          2389 => x"11",
          2390 => x"05",
          2391 => x"3f",
          2392 => x"08",
          2393 => x"da",
          2394 => x"71",
          2395 => x"84",
          2396 => x"3d",
          2397 => x"53",
          2398 => x"51",
          2399 => x"84",
          2400 => x"c6",
          2401 => x"39",
          2402 => x"80",
          2403 => x"7e",
          2404 => x"40",
          2405 => x"b8",
          2406 => x"11",
          2407 => x"05",
          2408 => x"3f",
          2409 => x"08",
          2410 => x"96",
          2411 => x"02",
          2412 => x"22",
          2413 => x"05",
          2414 => x"45",
          2415 => x"f0",
          2416 => x"80",
          2417 => x"bd",
          2418 => x"e4",
          2419 => x"38",
          2420 => x"b8",
          2421 => x"11",
          2422 => x"05",
          2423 => x"3f",
          2424 => x"08",
          2425 => x"dc",
          2426 => x"02",
          2427 => x"33",
          2428 => x"81",
          2429 => x"9b",
          2430 => x"fe",
          2431 => x"ff",
          2432 => x"e1",
          2433 => x"b8",
          2434 => x"2e",
          2435 => x"64",
          2436 => x"5d",
          2437 => x"70",
          2438 => x"e1",
          2439 => x"2e",
          2440 => x"f3",
          2441 => x"55",
          2442 => x"54",
          2443 => x"d7",
          2444 => x"51",
          2445 => x"f3",
          2446 => x"52",
          2447 => x"8a",
          2448 => x"39",
          2449 => x"51",
          2450 => x"f0",
          2451 => x"3d",
          2452 => x"53",
          2453 => x"51",
          2454 => x"84",
          2455 => x"80",
          2456 => x"64",
          2457 => x"ce",
          2458 => x"70",
          2459 => x"23",
          2460 => x"e7",
          2461 => x"e9",
          2462 => x"80",
          2463 => x"38",
          2464 => x"08",
          2465 => x"39",
          2466 => x"33",
          2467 => x"2e",
          2468 => x"f1",
          2469 => x"fc",
          2470 => x"d8",
          2471 => x"d6",
          2472 => x"f7",
          2473 => x"d8",
          2474 => x"ca",
          2475 => x"f6",
          2476 => x"f1",
          2477 => x"78",
          2478 => x"38",
          2479 => x"08",
          2480 => x"39",
          2481 => x"51",
          2482 => x"f9",
          2483 => x"f1",
          2484 => x"78",
          2485 => x"38",
          2486 => x"08",
          2487 => x"39",
          2488 => x"33",
          2489 => x"2e",
          2490 => x"f1",
          2491 => x"fb",
          2492 => x"f1",
          2493 => x"7d",
          2494 => x"38",
          2495 => x"08",
          2496 => x"39",
          2497 => x"33",
          2498 => x"2e",
          2499 => x"f1",
          2500 => x"fb",
          2501 => x"f1",
          2502 => x"7c",
          2503 => x"38",
          2504 => x"08",
          2505 => x"39",
          2506 => x"08",
          2507 => x"49",
          2508 => x"83",
          2509 => x"88",
          2510 => x"b5",
          2511 => x"0d",
          2512 => x"b9",
          2513 => x"c0",
          2514 => x"08",
          2515 => x"84",
          2516 => x"51",
          2517 => x"84",
          2518 => x"90",
          2519 => x"57",
          2520 => x"80",
          2521 => x"da",
          2522 => x"84",
          2523 => x"07",
          2524 => x"c0",
          2525 => x"08",
          2526 => x"84",
          2527 => x"51",
          2528 => x"84",
          2529 => x"90",
          2530 => x"57",
          2531 => x"80",
          2532 => x"da",
          2533 => x"84",
          2534 => x"07",
          2535 => x"80",
          2536 => x"c0",
          2537 => x"8c",
          2538 => x"87",
          2539 => x"0c",
          2540 => x"5c",
          2541 => x"5d",
          2542 => x"05",
          2543 => x"80",
          2544 => x"c4",
          2545 => x"70",
          2546 => x"70",
          2547 => x"d4",
          2548 => x"b6",
          2549 => x"83",
          2550 => x"3f",
          2551 => x"94",
          2552 => x"d2",
          2553 => x"d2",
          2554 => x"9f",
          2555 => x"d4",
          2556 => x"55",
          2557 => x"83",
          2558 => x"83",
          2559 => x"81",
          2560 => x"83",
          2561 => x"c4",
          2562 => x"97",
          2563 => x"3f",
          2564 => x"3d",
          2565 => x"08",
          2566 => x"75",
          2567 => x"73",
          2568 => x"38",
          2569 => x"81",
          2570 => x"52",
          2571 => x"09",
          2572 => x"38",
          2573 => x"33",
          2574 => x"06",
          2575 => x"70",
          2576 => x"38",
          2577 => x"06",
          2578 => x"2e",
          2579 => x"74",
          2580 => x"2e",
          2581 => x"80",
          2582 => x"81",
          2583 => x"54",
          2584 => x"2e",
          2585 => x"54",
          2586 => x"8b",
          2587 => x"2e",
          2588 => x"12",
          2589 => x"80",
          2590 => x"06",
          2591 => x"a0",
          2592 => x"06",
          2593 => x"54",
          2594 => x"70",
          2595 => x"25",
          2596 => x"52",
          2597 => x"2e",
          2598 => x"72",
          2599 => x"54",
          2600 => x"0c",
          2601 => x"84",
          2602 => x"87",
          2603 => x"70",
          2604 => x"38",
          2605 => x"ff",
          2606 => x"12",
          2607 => x"33",
          2608 => x"06",
          2609 => x"70",
          2610 => x"38",
          2611 => x"39",
          2612 => x"81",
          2613 => x"72",
          2614 => x"81",
          2615 => x"38",
          2616 => x"3d",
          2617 => x"72",
          2618 => x"80",
          2619 => x"e4",
          2620 => x"0d",
          2621 => x"fc",
          2622 => x"51",
          2623 => x"84",
          2624 => x"80",
          2625 => x"74",
          2626 => x"0c",
          2627 => x"04",
          2628 => x"76",
          2629 => x"ff",
          2630 => x"81",
          2631 => x"26",
          2632 => x"83",
          2633 => x"05",
          2634 => x"73",
          2635 => x"8a",
          2636 => x"33",
          2637 => x"70",
          2638 => x"fe",
          2639 => x"33",
          2640 => x"73",
          2641 => x"f2",
          2642 => x"33",
          2643 => x"74",
          2644 => x"e6",
          2645 => x"22",
          2646 => x"74",
          2647 => x"80",
          2648 => x"13",
          2649 => x"52",
          2650 => x"26",
          2651 => x"81",
          2652 => x"98",
          2653 => x"22",
          2654 => x"bc",
          2655 => x"33",
          2656 => x"b8",
          2657 => x"33",
          2658 => x"b4",
          2659 => x"33",
          2660 => x"b0",
          2661 => x"33",
          2662 => x"ac",
          2663 => x"33",
          2664 => x"a8",
          2665 => x"c0",
          2666 => x"73",
          2667 => x"a0",
          2668 => x"87",
          2669 => x"0c",
          2670 => x"84",
          2671 => x"86",
          2672 => x"f3",
          2673 => x"5b",
          2674 => x"9c",
          2675 => x"0c",
          2676 => x"bc",
          2677 => x"7b",
          2678 => x"98",
          2679 => x"7b",
          2680 => x"87",
          2681 => x"08",
          2682 => x"1c",
          2683 => x"98",
          2684 => x"7b",
          2685 => x"87",
          2686 => x"08",
          2687 => x"1c",
          2688 => x"98",
          2689 => x"7b",
          2690 => x"87",
          2691 => x"08",
          2692 => x"1c",
          2693 => x"98",
          2694 => x"79",
          2695 => x"80",
          2696 => x"83",
          2697 => x"59",
          2698 => x"ff",
          2699 => x"1b",
          2700 => x"1b",
          2701 => x"1b",
          2702 => x"1b",
          2703 => x"1b",
          2704 => x"83",
          2705 => x"52",
          2706 => x"51",
          2707 => x"3f",
          2708 => x"04",
          2709 => x"02",
          2710 => x"53",
          2711 => x"a8",
          2712 => x"80",
          2713 => x"84",
          2714 => x"98",
          2715 => x"2c",
          2716 => x"ff",
          2717 => x"06",
          2718 => x"83",
          2719 => x"71",
          2720 => x"0c",
          2721 => x"04",
          2722 => x"e8",
          2723 => x"b8",
          2724 => x"2b",
          2725 => x"51",
          2726 => x"2e",
          2727 => x"df",
          2728 => x"80",
          2729 => x"84",
          2730 => x"98",
          2731 => x"2c",
          2732 => x"ff",
          2733 => x"c7",
          2734 => x"0d",
          2735 => x"52",
          2736 => x"54",
          2737 => x"e7",
          2738 => x"b8",
          2739 => x"2b",
          2740 => x"51",
          2741 => x"2e",
          2742 => x"72",
          2743 => x"54",
          2744 => x"25",
          2745 => x"84",
          2746 => x"85",
          2747 => x"fc",
          2748 => x"9b",
          2749 => x"f1",
          2750 => x"81",
          2751 => x"55",
          2752 => x"2e",
          2753 => x"87",
          2754 => x"08",
          2755 => x"70",
          2756 => x"54",
          2757 => x"2e",
          2758 => x"91",
          2759 => x"06",
          2760 => x"e3",
          2761 => x"32",
          2762 => x"72",
          2763 => x"38",
          2764 => x"81",
          2765 => x"cf",
          2766 => x"ff",
          2767 => x"c0",
          2768 => x"70",
          2769 => x"38",
          2770 => x"90",
          2771 => x"0c",
          2772 => x"e4",
          2773 => x"0d",
          2774 => x"2a",
          2775 => x"51",
          2776 => x"38",
          2777 => x"81",
          2778 => x"80",
          2779 => x"71",
          2780 => x"06",
          2781 => x"2e",
          2782 => x"c0",
          2783 => x"70",
          2784 => x"81",
          2785 => x"52",
          2786 => x"d8",
          2787 => x"0d",
          2788 => x"33",
          2789 => x"9f",
          2790 => x"52",
          2791 => x"9c",
          2792 => x"0d",
          2793 => x"0d",
          2794 => x"75",
          2795 => x"52",
          2796 => x"2e",
          2797 => x"81",
          2798 => x"9c",
          2799 => x"ff",
          2800 => x"55",
          2801 => x"80",
          2802 => x"c0",
          2803 => x"70",
          2804 => x"81",
          2805 => x"52",
          2806 => x"8c",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"38",
          2810 => x"81",
          2811 => x"80",
          2812 => x"71",
          2813 => x"06",
          2814 => x"38",
          2815 => x"06",
          2816 => x"94",
          2817 => x"80",
          2818 => x"87",
          2819 => x"52",
          2820 => x"81",
          2821 => x"55",
          2822 => x"9b",
          2823 => x"b8",
          2824 => x"3d",
          2825 => x"91",
          2826 => x"06",
          2827 => x"98",
          2828 => x"32",
          2829 => x"72",
          2830 => x"38",
          2831 => x"81",
          2832 => x"80",
          2833 => x"38",
          2834 => x"84",
          2835 => x"2a",
          2836 => x"53",
          2837 => x"ce",
          2838 => x"ff",
          2839 => x"c0",
          2840 => x"70",
          2841 => x"06",
          2842 => x"80",
          2843 => x"38",
          2844 => x"a4",
          2845 => x"a0",
          2846 => x"9e",
          2847 => x"f1",
          2848 => x"c0",
          2849 => x"83",
          2850 => x"87",
          2851 => x"08",
          2852 => x"0c",
          2853 => x"9c",
          2854 => x"b0",
          2855 => x"9e",
          2856 => x"f1",
          2857 => x"c0",
          2858 => x"83",
          2859 => x"87",
          2860 => x"08",
          2861 => x"0c",
          2862 => x"b4",
          2863 => x"c0",
          2864 => x"9e",
          2865 => x"f1",
          2866 => x"c0",
          2867 => x"83",
          2868 => x"87",
          2869 => x"08",
          2870 => x"0c",
          2871 => x"c4",
          2872 => x"d0",
          2873 => x"9e",
          2874 => x"71",
          2875 => x"23",
          2876 => x"84",
          2877 => x"d8",
          2878 => x"9e",
          2879 => x"f1",
          2880 => x"c0",
          2881 => x"83",
          2882 => x"81",
          2883 => x"e4",
          2884 => x"87",
          2885 => x"08",
          2886 => x"0a",
          2887 => x"52",
          2888 => x"38",
          2889 => x"e5",
          2890 => x"87",
          2891 => x"08",
          2892 => x"0a",
          2893 => x"52",
          2894 => x"83",
          2895 => x"71",
          2896 => x"34",
          2897 => x"c0",
          2898 => x"70",
          2899 => x"06",
          2900 => x"70",
          2901 => x"38",
          2902 => x"83",
          2903 => x"80",
          2904 => x"9e",
          2905 => x"88",
          2906 => x"51",
          2907 => x"80",
          2908 => x"81",
          2909 => x"f1",
          2910 => x"0b",
          2911 => x"90",
          2912 => x"80",
          2913 => x"52",
          2914 => x"2e",
          2915 => x"52",
          2916 => x"e9",
          2917 => x"87",
          2918 => x"08",
          2919 => x"80",
          2920 => x"52",
          2921 => x"83",
          2922 => x"71",
          2923 => x"34",
          2924 => x"c0",
          2925 => x"70",
          2926 => x"06",
          2927 => x"70",
          2928 => x"38",
          2929 => x"83",
          2930 => x"80",
          2931 => x"9e",
          2932 => x"82",
          2933 => x"51",
          2934 => x"80",
          2935 => x"81",
          2936 => x"f1",
          2937 => x"0b",
          2938 => x"90",
          2939 => x"80",
          2940 => x"52",
          2941 => x"2e",
          2942 => x"52",
          2943 => x"ed",
          2944 => x"87",
          2945 => x"08",
          2946 => x"80",
          2947 => x"52",
          2948 => x"83",
          2949 => x"71",
          2950 => x"34",
          2951 => x"c0",
          2952 => x"70",
          2953 => x"51",
          2954 => x"80",
          2955 => x"81",
          2956 => x"f1",
          2957 => x"c0",
          2958 => x"98",
          2959 => x"8a",
          2960 => x"71",
          2961 => x"34",
          2962 => x"c0",
          2963 => x"70",
          2964 => x"51",
          2965 => x"80",
          2966 => x"81",
          2967 => x"f1",
          2968 => x"c0",
          2969 => x"83",
          2970 => x"84",
          2971 => x"71",
          2972 => x"34",
          2973 => x"c0",
          2974 => x"70",
          2975 => x"52",
          2976 => x"2e",
          2977 => x"52",
          2978 => x"f3",
          2979 => x"9e",
          2980 => x"06",
          2981 => x"f1",
          2982 => x"3d",
          2983 => x"52",
          2984 => x"fb",
          2985 => x"d8",
          2986 => x"b6",
          2987 => x"f1",
          2988 => x"73",
          2989 => x"83",
          2990 => x"c3",
          2991 => x"f1",
          2992 => x"74",
          2993 => x"83",
          2994 => x"54",
          2995 => x"38",
          2996 => x"33",
          2997 => x"a8",
          2998 => x"e9",
          2999 => x"84",
          3000 => x"f1",
          3001 => x"73",
          3002 => x"83",
          3003 => x"56",
          3004 => x"38",
          3005 => x"33",
          3006 => x"90",
          3007 => x"f1",
          3008 => x"83",
          3009 => x"f1",
          3010 => x"75",
          3011 => x"83",
          3012 => x"54",
          3013 => x"38",
          3014 => x"33",
          3015 => x"93",
          3016 => x"ed",
          3017 => x"82",
          3018 => x"f1",
          3019 => x"73",
          3020 => x"83",
          3021 => x"c2",
          3022 => x"f1",
          3023 => x"83",
          3024 => x"ff",
          3025 => x"83",
          3026 => x"52",
          3027 => x"51",
          3028 => x"3f",
          3029 => x"08",
          3030 => x"a8",
          3031 => x"ab",
          3032 => x"d0",
          3033 => x"3f",
          3034 => x"22",
          3035 => x"d8",
          3036 => x"97",
          3037 => x"d8",
          3038 => x"84",
          3039 => x"51",
          3040 => x"84",
          3041 => x"bd",
          3042 => x"76",
          3043 => x"54",
          3044 => x"08",
          3045 => x"80",
          3046 => x"ef",
          3047 => x"eb",
          3048 => x"80",
          3049 => x"f1",
          3050 => x"74",
          3051 => x"51",
          3052 => x"87",
          3053 => x"83",
          3054 => x"56",
          3055 => x"52",
          3056 => x"e4",
          3057 => x"e4",
          3058 => x"c0",
          3059 => x"31",
          3060 => x"b8",
          3061 => x"83",
          3062 => x"ff",
          3063 => x"8a",
          3064 => x"3f",
          3065 => x"04",
          3066 => x"08",
          3067 => x"c0",
          3068 => x"c9",
          3069 => x"b8",
          3070 => x"84",
          3071 => x"71",
          3072 => x"84",
          3073 => x"52",
          3074 => x"51",
          3075 => x"3f",
          3076 => x"33",
          3077 => x"2e",
          3078 => x"ff",
          3079 => x"db",
          3080 => x"d2",
          3081 => x"cc",
          3082 => x"3f",
          3083 => x"08",
          3084 => x"d8",
          3085 => x"d3",
          3086 => x"cc",
          3087 => x"d9",
          3088 => x"b3",
          3089 => x"f1",
          3090 => x"83",
          3091 => x"ff",
          3092 => x"83",
          3093 => x"c0",
          3094 => x"f1",
          3095 => x"83",
          3096 => x"ff",
          3097 => x"83",
          3098 => x"56",
          3099 => x"52",
          3100 => x"b4",
          3101 => x"e4",
          3102 => x"c0",
          3103 => x"31",
          3104 => x"b8",
          3105 => x"83",
          3106 => x"ff",
          3107 => x"83",
          3108 => x"55",
          3109 => x"fe",
          3110 => x"cc",
          3111 => x"8c",
          3112 => x"d2",
          3113 => x"ee",
          3114 => x"80",
          3115 => x"38",
          3116 => x"83",
          3117 => x"ff",
          3118 => x"83",
          3119 => x"56",
          3120 => x"fc",
          3121 => x"39",
          3122 => x"51",
          3123 => x"3f",
          3124 => x"33",
          3125 => x"2e",
          3126 => x"d7",
          3127 => x"ac",
          3128 => x"92",
          3129 => x"e7",
          3130 => x"80",
          3131 => x"38",
          3132 => x"f1",
          3133 => x"83",
          3134 => x"ff",
          3135 => x"83",
          3136 => x"56",
          3137 => x"fc",
          3138 => x"39",
          3139 => x"33",
          3140 => x"e0",
          3141 => x"f3",
          3142 => x"f1",
          3143 => x"80",
          3144 => x"38",
          3145 => x"f1",
          3146 => x"83",
          3147 => x"ff",
          3148 => x"83",
          3149 => x"54",
          3150 => x"fb",
          3151 => x"39",
          3152 => x"08",
          3153 => x"08",
          3154 => x"83",
          3155 => x"ff",
          3156 => x"83",
          3157 => x"56",
          3158 => x"fb",
          3159 => x"39",
          3160 => x"08",
          3161 => x"08",
          3162 => x"83",
          3163 => x"ff",
          3164 => x"83",
          3165 => x"54",
          3166 => x"fa",
          3167 => x"39",
          3168 => x"08",
          3169 => x"08",
          3170 => x"83",
          3171 => x"ff",
          3172 => x"83",
          3173 => x"55",
          3174 => x"fa",
          3175 => x"39",
          3176 => x"08",
          3177 => x"08",
          3178 => x"83",
          3179 => x"ff",
          3180 => x"83",
          3181 => x"56",
          3182 => x"fa",
          3183 => x"39",
          3184 => x"08",
          3185 => x"08",
          3186 => x"83",
          3187 => x"ff",
          3188 => x"83",
          3189 => x"54",
          3190 => x"f9",
          3191 => x"39",
          3192 => x"51",
          3193 => x"3f",
          3194 => x"51",
          3195 => x"3f",
          3196 => x"33",
          3197 => x"2e",
          3198 => x"c4",
          3199 => x"0d",
          3200 => x"33",
          3201 => x"26",
          3202 => x"10",
          3203 => x"ec",
          3204 => x"08",
          3205 => x"c0",
          3206 => x"ef",
          3207 => x"0d",
          3208 => x"c8",
          3209 => x"e3",
          3210 => x"0d",
          3211 => x"d0",
          3212 => x"d7",
          3213 => x"0d",
          3214 => x"d8",
          3215 => x"cb",
          3216 => x"0d",
          3217 => x"e0",
          3218 => x"bf",
          3219 => x"0d",
          3220 => x"e8",
          3221 => x"b3",
          3222 => x"0d",
          3223 => x"80",
          3224 => x"0b",
          3225 => x"84",
          3226 => x"f1",
          3227 => x"c0",
          3228 => x"04",
          3229 => x"aa",
          3230 => x"3d",
          3231 => x"81",
          3232 => x"80",
          3233 => x"d0",
          3234 => x"88",
          3235 => x"b8",
          3236 => x"ed",
          3237 => x"57",
          3238 => x"f2",
          3239 => x"55",
          3240 => x"76",
          3241 => x"8f",
          3242 => x"e4",
          3243 => x"a4",
          3244 => x"c0",
          3245 => x"b8",
          3246 => x"17",
          3247 => x"0b",
          3248 => x"08",
          3249 => x"84",
          3250 => x"ff",
          3251 => x"55",
          3252 => x"34",
          3253 => x"30",
          3254 => x"9f",
          3255 => x"55",
          3256 => x"85",
          3257 => x"b0",
          3258 => x"d0",
          3259 => x"08",
          3260 => x"87",
          3261 => x"b8",
          3262 => x"38",
          3263 => x"9a",
          3264 => x"b8",
          3265 => x"3d",
          3266 => x"e1",
          3267 => x"ad",
          3268 => x"76",
          3269 => x"06",
          3270 => x"52",
          3271 => x"aa",
          3272 => x"c0",
          3273 => x"3d",
          3274 => x"b8",
          3275 => x"34",
          3276 => x"e1",
          3277 => x"ad",
          3278 => x"0b",
          3279 => x"0c",
          3280 => x"04",
          3281 => x"ab",
          3282 => x"3d",
          3283 => x"5d",
          3284 => x"57",
          3285 => x"a0",
          3286 => x"38",
          3287 => x"3d",
          3288 => x"10",
          3289 => x"f2",
          3290 => x"08",
          3291 => x"bf",
          3292 => x"b8",
          3293 => x"79",
          3294 => x"51",
          3295 => x"84",
          3296 => x"90",
          3297 => x"33",
          3298 => x"2e",
          3299 => x"73",
          3300 => x"38",
          3301 => x"81",
          3302 => x"54",
          3303 => x"c2",
          3304 => x"73",
          3305 => x"0c",
          3306 => x"04",
          3307 => x"aa",
          3308 => x"11",
          3309 => x"05",
          3310 => x"3f",
          3311 => x"08",
          3312 => x"38",
          3313 => x"78",
          3314 => x"fd",
          3315 => x"b8",
          3316 => x"ff",
          3317 => x"80",
          3318 => x"81",
          3319 => x"ff",
          3320 => x"82",
          3321 => x"fa",
          3322 => x"39",
          3323 => x"05",
          3324 => x"27",
          3325 => x"81",
          3326 => x"70",
          3327 => x"73",
          3328 => x"81",
          3329 => x"38",
          3330 => x"eb",
          3331 => x"8d",
          3332 => x"fe",
          3333 => x"84",
          3334 => x"53",
          3335 => x"08",
          3336 => x"84",
          3337 => x"b8",
          3338 => x"d0",
          3339 => x"d0",
          3340 => x"f8",
          3341 => x"82",
          3342 => x"84",
          3343 => x"80",
          3344 => x"77",
          3345 => x"e3",
          3346 => x"e4",
          3347 => x"0b",
          3348 => x"08",
          3349 => x"84",
          3350 => x"ff",
          3351 => x"58",
          3352 => x"34",
          3353 => x"52",
          3354 => x"e1",
          3355 => x"ff",
          3356 => x"74",
          3357 => x"81",
          3358 => x"38",
          3359 => x"b8",
          3360 => x"3d",
          3361 => x"3d",
          3362 => x"08",
          3363 => x"b9",
          3364 => x"41",
          3365 => x"b4",
          3366 => x"f2",
          3367 => x"f2",
          3368 => x"5d",
          3369 => x"74",
          3370 => x"33",
          3371 => x"80",
          3372 => x"38",
          3373 => x"91",
          3374 => x"70",
          3375 => x"57",
          3376 => x"38",
          3377 => x"90",
          3378 => x"3d",
          3379 => x"5f",
          3380 => x"80",
          3381 => x"e4",
          3382 => x"70",
          3383 => x"56",
          3384 => x"ec",
          3385 => x"ff",
          3386 => x"a0",
          3387 => x"2b",
          3388 => x"84",
          3389 => x"70",
          3390 => x"97",
          3391 => x"2c",
          3392 => x"10",
          3393 => x"05",
          3394 => x"70",
          3395 => x"5c",
          3396 => x"5b",
          3397 => x"81",
          3398 => x"2e",
          3399 => x"78",
          3400 => x"87",
          3401 => x"80",
          3402 => x"ff",
          3403 => x"98",
          3404 => x"80",
          3405 => x"cb",
          3406 => x"16",
          3407 => x"56",
          3408 => x"83",
          3409 => x"33",
          3410 => x"61",
          3411 => x"83",
          3412 => x"08",
          3413 => x"56",
          3414 => x"2e",
          3415 => x"76",
          3416 => x"38",
          3417 => x"9c",
          3418 => x"76",
          3419 => x"99",
          3420 => x"70",
          3421 => x"98",
          3422 => x"9c",
          3423 => x"2b",
          3424 => x"71",
          3425 => x"70",
          3426 => x"dd",
          3427 => x"5f",
          3428 => x"58",
          3429 => x"7a",
          3430 => x"90",
          3431 => x"d0",
          3432 => x"ac",
          3433 => x"76",
          3434 => x"75",
          3435 => x"29",
          3436 => x"05",
          3437 => x"70",
          3438 => x"59",
          3439 => x"95",
          3440 => x"38",
          3441 => x"70",
          3442 => x"55",
          3443 => x"dd",
          3444 => x"42",
          3445 => x"25",
          3446 => x"dd",
          3447 => x"18",
          3448 => x"55",
          3449 => x"ff",
          3450 => x"80",
          3451 => x"38",
          3452 => x"81",
          3453 => x"2e",
          3454 => x"fe",
          3455 => x"56",
          3456 => x"80",
          3457 => x"e9",
          3458 => x"d0",
          3459 => x"84",
          3460 => x"79",
          3461 => x"7f",
          3462 => x"74",
          3463 => x"b0",
          3464 => x"10",
          3465 => x"05",
          3466 => x"04",
          3467 => x"15",
          3468 => x"80",
          3469 => x"a0",
          3470 => x"84",
          3471 => x"d9",
          3472 => x"a8",
          3473 => x"80",
          3474 => x"38",
          3475 => x"08",
          3476 => x"ff",
          3477 => x"84",
          3478 => x"ff",
          3479 => x"84",
          3480 => x"fc",
          3481 => x"d0",
          3482 => x"81",
          3483 => x"d0",
          3484 => x"57",
          3485 => x"27",
          3486 => x"84",
          3487 => x"52",
          3488 => x"77",
          3489 => x"34",
          3490 => x"33",
          3491 => x"b5",
          3492 => x"bc",
          3493 => x"2e",
          3494 => x"7c",
          3495 => x"f2",
          3496 => x"08",
          3497 => x"8f",
          3498 => x"84",
          3499 => x"75",
          3500 => x"d0",
          3501 => x"d0",
          3502 => x"56",
          3503 => x"b6",
          3504 => x"c8",
          3505 => x"51",
          3506 => x"3f",
          3507 => x"08",
          3508 => x"ff",
          3509 => x"84",
          3510 => x"52",
          3511 => x"b5",
          3512 => x"d0",
          3513 => x"05",
          3514 => x"d0",
          3515 => x"81",
          3516 => x"74",
          3517 => x"51",
          3518 => x"3f",
          3519 => x"a8",
          3520 => x"39",
          3521 => x"83",
          3522 => x"56",
          3523 => x"38",
          3524 => x"83",
          3525 => x"fc",
          3526 => x"55",
          3527 => x"38",
          3528 => x"75",
          3529 => x"a8",
          3530 => x"ff",
          3531 => x"84",
          3532 => x"84",
          3533 => x"84",
          3534 => x"81",
          3535 => x"05",
          3536 => x"7b",
          3537 => x"a5",
          3538 => x"a4",
          3539 => x"a8",
          3540 => x"74",
          3541 => x"9e",
          3542 => x"c8",
          3543 => x"51",
          3544 => x"3f",
          3545 => x"08",
          3546 => x"ff",
          3547 => x"84",
          3548 => x"52",
          3549 => x"b3",
          3550 => x"d0",
          3551 => x"05",
          3552 => x"d0",
          3553 => x"81",
          3554 => x"c7",
          3555 => x"a8",
          3556 => x"ff",
          3557 => x"a4",
          3558 => x"55",
          3559 => x"fa",
          3560 => x"d4",
          3561 => x"81",
          3562 => x"84",
          3563 => x"7b",
          3564 => x"52",
          3565 => x"b9",
          3566 => x"a8",
          3567 => x"ff",
          3568 => x"a4",
          3569 => x"55",
          3570 => x"fa",
          3571 => x"d4",
          3572 => x"81",
          3573 => x"84",
          3574 => x"7b",
          3575 => x"52",
          3576 => x"8d",
          3577 => x"a8",
          3578 => x"ff",
          3579 => x"a4",
          3580 => x"55",
          3581 => x"ff",
          3582 => x"d4",
          3583 => x"a8",
          3584 => x"a4",
          3585 => x"74",
          3586 => x"c4",
          3587 => x"5b",
          3588 => x"a4",
          3589 => x"2b",
          3590 => x"7c",
          3591 => x"43",
          3592 => x"76",
          3593 => x"38",
          3594 => x"08",
          3595 => x"ff",
          3596 => x"84",
          3597 => x"70",
          3598 => x"98",
          3599 => x"a4",
          3600 => x"57",
          3601 => x"24",
          3602 => x"84",
          3603 => x"52",
          3604 => x"b2",
          3605 => x"81",
          3606 => x"81",
          3607 => x"70",
          3608 => x"d0",
          3609 => x"56",
          3610 => x"24",
          3611 => x"84",
          3612 => x"52",
          3613 => x"b1",
          3614 => x"81",
          3615 => x"81",
          3616 => x"70",
          3617 => x"d0",
          3618 => x"56",
          3619 => x"25",
          3620 => x"f8",
          3621 => x"16",
          3622 => x"33",
          3623 => x"d4",
          3624 => x"77",
          3625 => x"b1",
          3626 => x"81",
          3627 => x"81",
          3628 => x"70",
          3629 => x"d0",
          3630 => x"57",
          3631 => x"25",
          3632 => x"7b",
          3633 => x"18",
          3634 => x"84",
          3635 => x"52",
          3636 => x"ff",
          3637 => x"75",
          3638 => x"29",
          3639 => x"05",
          3640 => x"84",
          3641 => x"5b",
          3642 => x"76",
          3643 => x"38",
          3644 => x"84",
          3645 => x"55",
          3646 => x"f7",
          3647 => x"d4",
          3648 => x"88",
          3649 => x"e9",
          3650 => x"a8",
          3651 => x"57",
          3652 => x"a8",
          3653 => x"ff",
          3654 => x"39",
          3655 => x"33",
          3656 => x"80",
          3657 => x"d4",
          3658 => x"8a",
          3659 => x"c1",
          3660 => x"a4",
          3661 => x"f4",
          3662 => x"b8",
          3663 => x"ff",
          3664 => x"89",
          3665 => x"d0",
          3666 => x"76",
          3667 => x"d8",
          3668 => x"d4",
          3669 => x"10",
          3670 => x"05",
          3671 => x"5e",
          3672 => x"a0",
          3673 => x"2b",
          3674 => x"83",
          3675 => x"81",
          3676 => x"57",
          3677 => x"fb",
          3678 => x"e4",
          3679 => x"83",
          3680 => x"70",
          3681 => x"f1",
          3682 => x"08",
          3683 => x"74",
          3684 => x"83",
          3685 => x"56",
          3686 => x"8c",
          3687 => x"cc",
          3688 => x"80",
          3689 => x"38",
          3690 => x"d0",
          3691 => x"0b",
          3692 => x"34",
          3693 => x"e4",
          3694 => x"0d",
          3695 => x"a8",
          3696 => x"80",
          3697 => x"84",
          3698 => x"52",
          3699 => x"af",
          3700 => x"d4",
          3701 => x"a0",
          3702 => x"95",
          3703 => x"c8",
          3704 => x"51",
          3705 => x"3f",
          3706 => x"33",
          3707 => x"75",
          3708 => x"34",
          3709 => x"06",
          3710 => x"38",
          3711 => x"51",
          3712 => x"3f",
          3713 => x"d0",
          3714 => x"0b",
          3715 => x"34",
          3716 => x"83",
          3717 => x"0b",
          3718 => x"84",
          3719 => x"55",
          3720 => x"b6",
          3721 => x"c8",
          3722 => x"51",
          3723 => x"3f",
          3724 => x"08",
          3725 => x"ff",
          3726 => x"84",
          3727 => x"52",
          3728 => x"ae",
          3729 => x"d0",
          3730 => x"05",
          3731 => x"d0",
          3732 => x"81",
          3733 => x"74",
          3734 => x"d1",
          3735 => x"9f",
          3736 => x"0b",
          3737 => x"34",
          3738 => x"d0",
          3739 => x"84",
          3740 => x"b4",
          3741 => x"84",
          3742 => x"70",
          3743 => x"5c",
          3744 => x"2e",
          3745 => x"84",
          3746 => x"ff",
          3747 => x"84",
          3748 => x"ff",
          3749 => x"84",
          3750 => x"84",
          3751 => x"52",
          3752 => x"ad",
          3753 => x"d0",
          3754 => x"98",
          3755 => x"2c",
          3756 => x"33",
          3757 => x"56",
          3758 => x"80",
          3759 => x"d4",
          3760 => x"a0",
          3761 => x"a9",
          3762 => x"a8",
          3763 => x"2b",
          3764 => x"84",
          3765 => x"5d",
          3766 => x"74",
          3767 => x"f0",
          3768 => x"c8",
          3769 => x"51",
          3770 => x"3f",
          3771 => x"0a",
          3772 => x"0a",
          3773 => x"2c",
          3774 => x"33",
          3775 => x"74",
          3776 => x"cc",
          3777 => x"c8",
          3778 => x"51",
          3779 => x"3f",
          3780 => x"0a",
          3781 => x"0a",
          3782 => x"2c",
          3783 => x"33",
          3784 => x"78",
          3785 => x"b9",
          3786 => x"39",
          3787 => x"81",
          3788 => x"34",
          3789 => x"08",
          3790 => x"51",
          3791 => x"3f",
          3792 => x"0a",
          3793 => x"0a",
          3794 => x"2c",
          3795 => x"33",
          3796 => x"75",
          3797 => x"e6",
          3798 => x"57",
          3799 => x"77",
          3800 => x"c8",
          3801 => x"33",
          3802 => x"85",
          3803 => x"80",
          3804 => x"80",
          3805 => x"98",
          3806 => x"a4",
          3807 => x"5b",
          3808 => x"ff",
          3809 => x"b6",
          3810 => x"a8",
          3811 => x"ff",
          3812 => x"76",
          3813 => x"b8",
          3814 => x"a4",
          3815 => x"75",
          3816 => x"74",
          3817 => x"98",
          3818 => x"76",
          3819 => x"38",
          3820 => x"7a",
          3821 => x"34",
          3822 => x"0a",
          3823 => x"0a",
          3824 => x"2c",
          3825 => x"33",
          3826 => x"75",
          3827 => x"38",
          3828 => x"74",
          3829 => x"34",
          3830 => x"06",
          3831 => x"b3",
          3832 => x"34",
          3833 => x"33",
          3834 => x"25",
          3835 => x"17",
          3836 => x"d0",
          3837 => x"57",
          3838 => x"33",
          3839 => x"0a",
          3840 => x"0a",
          3841 => x"2c",
          3842 => x"06",
          3843 => x"58",
          3844 => x"81",
          3845 => x"98",
          3846 => x"2c",
          3847 => x"06",
          3848 => x"75",
          3849 => x"a8",
          3850 => x"c8",
          3851 => x"51",
          3852 => x"3f",
          3853 => x"0a",
          3854 => x"0a",
          3855 => x"2c",
          3856 => x"33",
          3857 => x"75",
          3858 => x"84",
          3859 => x"c8",
          3860 => x"51",
          3861 => x"3f",
          3862 => x"0a",
          3863 => x"0a",
          3864 => x"2c",
          3865 => x"33",
          3866 => x"74",
          3867 => x"b9",
          3868 => x"39",
          3869 => x"08",
          3870 => x"2e",
          3871 => x"75",
          3872 => x"a7",
          3873 => x"e4",
          3874 => x"a4",
          3875 => x"e4",
          3876 => x"06",
          3877 => x"75",
          3878 => x"ff",
          3879 => x"84",
          3880 => x"84",
          3881 => x"56",
          3882 => x"2e",
          3883 => x"84",
          3884 => x"52",
          3885 => x"a9",
          3886 => x"d4",
          3887 => x"a0",
          3888 => x"ad",
          3889 => x"c8",
          3890 => x"51",
          3891 => x"3f",
          3892 => x"33",
          3893 => x"7a",
          3894 => x"34",
          3895 => x"06",
          3896 => x"a8",
          3897 => x"8b",
          3898 => x"e4",
          3899 => x"d0",
          3900 => x"e4",
          3901 => x"38",
          3902 => x"cc",
          3903 => x"ca",
          3904 => x"39",
          3905 => x"08",
          3906 => x"70",
          3907 => x"ff",
          3908 => x"75",
          3909 => x"29",
          3910 => x"05",
          3911 => x"84",
          3912 => x"52",
          3913 => x"76",
          3914 => x"84",
          3915 => x"70",
          3916 => x"98",
          3917 => x"ff",
          3918 => x"5a",
          3919 => x"25",
          3920 => x"fd",
          3921 => x"f2",
          3922 => x"2e",
          3923 => x"83",
          3924 => x"93",
          3925 => x"55",
          3926 => x"ff",
          3927 => x"58",
          3928 => x"25",
          3929 => x"0b",
          3930 => x"34",
          3931 => x"08",
          3932 => x"2e",
          3933 => x"74",
          3934 => x"f6",
          3935 => x"d0",
          3936 => x"d9",
          3937 => x"0b",
          3938 => x"0c",
          3939 => x"3d",
          3940 => x"bc",
          3941 => x"80",
          3942 => x"80",
          3943 => x"16",
          3944 => x"56",
          3945 => x"ff",
          3946 => x"ba",
          3947 => x"ff",
          3948 => x"84",
          3949 => x"84",
          3950 => x"84",
          3951 => x"81",
          3952 => x"05",
          3953 => x"7b",
          3954 => x"a1",
          3955 => x"84",
          3956 => x"84",
          3957 => x"57",
          3958 => x"80",
          3959 => x"38",
          3960 => x"08",
          3961 => x"ff",
          3962 => x"84",
          3963 => x"52",
          3964 => x"a6",
          3965 => x"d4",
          3966 => x"88",
          3967 => x"f1",
          3968 => x"a8",
          3969 => x"5a",
          3970 => x"a8",
          3971 => x"ff",
          3972 => x"39",
          3973 => x"80",
          3974 => x"a8",
          3975 => x"84",
          3976 => x"7b",
          3977 => x"0c",
          3978 => x"04",
          3979 => x"a9",
          3980 => x"b8",
          3981 => x"d0",
          3982 => x"b8",
          3983 => x"ff",
          3984 => x"53",
          3985 => x"51",
          3986 => x"3f",
          3987 => x"81",
          3988 => x"d0",
          3989 => x"d0",
          3990 => x"52",
          3991 => x"80",
          3992 => x"38",
          3993 => x"08",
          3994 => x"ff",
          3995 => x"84",
          3996 => x"52",
          3997 => x"a5",
          3998 => x"d4",
          3999 => x"88",
          4000 => x"ed",
          4001 => x"a8",
          4002 => x"57",
          4003 => x"a8",
          4004 => x"ff",
          4005 => x"39",
          4006 => x"a9",
          4007 => x"b8",
          4008 => x"d0",
          4009 => x"b8",
          4010 => x"ff",
          4011 => x"53",
          4012 => x"51",
          4013 => x"3f",
          4014 => x"81",
          4015 => x"d0",
          4016 => x"d0",
          4017 => x"58",
          4018 => x"80",
          4019 => x"38",
          4020 => x"08",
          4021 => x"ff",
          4022 => x"84",
          4023 => x"52",
          4024 => x"a5",
          4025 => x"d4",
          4026 => x"88",
          4027 => x"81",
          4028 => x"a8",
          4029 => x"41",
          4030 => x"a8",
          4031 => x"ff",
          4032 => x"39",
          4033 => x"d6",
          4034 => x"f2",
          4035 => x"82",
          4036 => x"06",
          4037 => x"05",
          4038 => x"54",
          4039 => x"80",
          4040 => x"84",
          4041 => x"7b",
          4042 => x"d4",
          4043 => x"10",
          4044 => x"05",
          4045 => x"41",
          4046 => x"2e",
          4047 => x"75",
          4048 => x"74",
          4049 => x"a5",
          4050 => x"d4",
          4051 => x"70",
          4052 => x"5a",
          4053 => x"27",
          4054 => x"77",
          4055 => x"34",
          4056 => x"b4",
          4057 => x"05",
          4058 => x"7b",
          4059 => x"81",
          4060 => x"83",
          4061 => x"52",
          4062 => x"ba",
          4063 => x"f2",
          4064 => x"81",
          4065 => x"80",
          4066 => x"a8",
          4067 => x"84",
          4068 => x"7b",
          4069 => x"0c",
          4070 => x"04",
          4071 => x"52",
          4072 => x"08",
          4073 => x"f8",
          4074 => x"e4",
          4075 => x"38",
          4076 => x"08",
          4077 => x"5d",
          4078 => x"08",
          4079 => x"52",
          4080 => x"b7",
          4081 => x"b8",
          4082 => x"84",
          4083 => x"7b",
          4084 => x"06",
          4085 => x"84",
          4086 => x"51",
          4087 => x"3f",
          4088 => x"08",
          4089 => x"84",
          4090 => x"25",
          4091 => x"84",
          4092 => x"ff",
          4093 => x"58",
          4094 => x"34",
          4095 => x"06",
          4096 => x"33",
          4097 => x"83",
          4098 => x"70",
          4099 => x"58",
          4100 => x"f2",
          4101 => x"2b",
          4102 => x"83",
          4103 => x"81",
          4104 => x"58",
          4105 => x"cb",
          4106 => x"e4",
          4107 => x"83",
          4108 => x"70",
          4109 => x"f1",
          4110 => x"08",
          4111 => x"74",
          4112 => x"1d",
          4113 => x"06",
          4114 => x"7d",
          4115 => x"80",
          4116 => x"2e",
          4117 => x"fe",
          4118 => x"e8",
          4119 => x"e6",
          4120 => x"79",
          4121 => x"ff",
          4122 => x"83",
          4123 => x"81",
          4124 => x"ff",
          4125 => x"93",
          4126 => x"c8",
          4127 => x"83",
          4128 => x"ff",
          4129 => x"51",
          4130 => x"3f",
          4131 => x"33",
          4132 => x"87",
          4133 => x"f1",
          4134 => x"1b",
          4135 => x"56",
          4136 => x"cf",
          4137 => x"e4",
          4138 => x"83",
          4139 => x"70",
          4140 => x"f1",
          4141 => x"08",
          4142 => x"74",
          4143 => x"82",
          4144 => x"39",
          4145 => x"d4",
          4146 => x"39",
          4147 => x"d4",
          4148 => x"39",
          4149 => x"51",
          4150 => x"3f",
          4151 => x"38",
          4152 => x"f2",
          4153 => x"80",
          4154 => x"02",
          4155 => x"c7",
          4156 => x"53",
          4157 => x"81",
          4158 => x"81",
          4159 => x"38",
          4160 => x"83",
          4161 => x"82",
          4162 => x"38",
          4163 => x"80",
          4164 => x"b0",
          4165 => x"57",
          4166 => x"a0",
          4167 => x"2e",
          4168 => x"83",
          4169 => x"75",
          4170 => x"34",
          4171 => x"92",
          4172 => x"90",
          4173 => x"2b",
          4174 => x"07",
          4175 => x"07",
          4176 => x"7f",
          4177 => x"5b",
          4178 => x"94",
          4179 => x"70",
          4180 => x"0c",
          4181 => x"84",
          4182 => x"76",
          4183 => x"38",
          4184 => x"a2",
          4185 => x"90",
          4186 => x"b6",
          4187 => x"31",
          4188 => x"a0",
          4189 => x"15",
          4190 => x"70",
          4191 => x"34",
          4192 => x"72",
          4193 => x"3d",
          4194 => x"a7",
          4195 => x"83",
          4196 => x"70",
          4197 => x"83",
          4198 => x"71",
          4199 => x"74",
          4200 => x"58",
          4201 => x"a7",
          4202 => x"84",
          4203 => x"70",
          4204 => x"84",
          4205 => x"70",
          4206 => x"83",
          4207 => x"70",
          4208 => x"06",
          4209 => x"5d",
          4210 => x"5e",
          4211 => x"73",
          4212 => x"38",
          4213 => x"75",
          4214 => x"81",
          4215 => x"81",
          4216 => x"81",
          4217 => x"83",
          4218 => x"62",
          4219 => x"70",
          4220 => x"5d",
          4221 => x"5b",
          4222 => x"26",
          4223 => x"f8",
          4224 => x"76",
          4225 => x"7d",
          4226 => x"5f",
          4227 => x"5c",
          4228 => x"fe",
          4229 => x"7d",
          4230 => x"77",
          4231 => x"38",
          4232 => x"81",
          4233 => x"83",
          4234 => x"74",
          4235 => x"56",
          4236 => x"86",
          4237 => x"59",
          4238 => x"80",
          4239 => x"d8",
          4240 => x"ff",
          4241 => x"d7",
          4242 => x"ff",
          4243 => x"92",
          4244 => x"29",
          4245 => x"57",
          4246 => x"57",
          4247 => x"81",
          4248 => x"81",
          4249 => x"81",
          4250 => x"71",
          4251 => x"54",
          4252 => x"2e",
          4253 => x"80",
          4254 => x"94",
          4255 => x"83",
          4256 => x"83",
          4257 => x"70",
          4258 => x"90",
          4259 => x"88",
          4260 => x"07",
          4261 => x"56",
          4262 => x"79",
          4263 => x"38",
          4264 => x"72",
          4265 => x"83",
          4266 => x"70",
          4267 => x"70",
          4268 => x"83",
          4269 => x"71",
          4270 => x"86",
          4271 => x"11",
          4272 => x"56",
          4273 => x"a7",
          4274 => x"14",
          4275 => x"33",
          4276 => x"06",
          4277 => x"33",
          4278 => x"06",
          4279 => x"22",
          4280 => x"ff",
          4281 => x"29",
          4282 => x"5a",
          4283 => x"5f",
          4284 => x"79",
          4285 => x"38",
          4286 => x"15",
          4287 => x"19",
          4288 => x"81",
          4289 => x"81",
          4290 => x"71",
          4291 => x"ff",
          4292 => x"81",
          4293 => x"75",
          4294 => x"5b",
          4295 => x"7b",
          4296 => x"38",
          4297 => x"53",
          4298 => x"16",
          4299 => x"5b",
          4300 => x"e2",
          4301 => x"06",
          4302 => x"da",
          4303 => x"39",
          4304 => x"7b",
          4305 => x"9a",
          4306 => x"0d",
          4307 => x"8c",
          4308 => x"73",
          4309 => x"34",
          4310 => x"81",
          4311 => x"ee",
          4312 => x"80",
          4313 => x"ff",
          4314 => x"86",
          4315 => x"56",
          4316 => x"80",
          4317 => x"ee",
          4318 => x"8a",
          4319 => x"74",
          4320 => x"75",
          4321 => x"83",
          4322 => x"3f",
          4323 => x"e0",
          4324 => x"54",
          4325 => x"86",
          4326 => x"73",
          4327 => x"07",
          4328 => x"75",
          4329 => x"70",
          4330 => x"80",
          4331 => x"53",
          4332 => x"86",
          4333 => x"08",
          4334 => x"81",
          4335 => x"72",
          4336 => x"f3",
          4337 => x"81",
          4338 => x"07",
          4339 => x"34",
          4340 => x"84",
          4341 => x"80",
          4342 => x"e4",
          4343 => x"0d",
          4344 => x"d8",
          4345 => x"e4",
          4346 => x"3d",
          4347 => x"05",
          4348 => x"05",
          4349 => x"84",
          4350 => x"5b",
          4351 => x"53",
          4352 => x"82",
          4353 => x"b6",
          4354 => x"f8",
          4355 => x"f8",
          4356 => x"71",
          4357 => x"a7",
          4358 => x"83",
          4359 => x"5f",
          4360 => x"71",
          4361 => x"70",
          4362 => x"06",
          4363 => x"33",
          4364 => x"53",
          4365 => x"83",
          4366 => x"f8",
          4367 => x"05",
          4368 => x"f8",
          4369 => x"f8",
          4370 => x"05",
          4371 => x"06",
          4372 => x"06",
          4373 => x"72",
          4374 => x"8c",
          4375 => x"53",
          4376 => x"94",
          4377 => x"92",
          4378 => x"ff",
          4379 => x"b6",
          4380 => x"55",
          4381 => x"26",
          4382 => x"84",
          4383 => x"76",
          4384 => x"58",
          4385 => x"9f",
          4386 => x"38",
          4387 => x"70",
          4388 => x"e0",
          4389 => x"e0",
          4390 => x"72",
          4391 => x"54",
          4392 => x"81",
          4393 => x"81",
          4394 => x"b6",
          4395 => x"e3",
          4396 => x"9f",
          4397 => x"83",
          4398 => x"84",
          4399 => x"54",
          4400 => x"e0",
          4401 => x"74",
          4402 => x"05",
          4403 => x"14",
          4404 => x"74",
          4405 => x"84",
          4406 => x"ff",
          4407 => x"83",
          4408 => x"75",
          4409 => x"ff",
          4410 => x"ff",
          4411 => x"54",
          4412 => x"81",
          4413 => x"74",
          4414 => x"84",
          4415 => x"71",
          4416 => x"55",
          4417 => x"86",
          4418 => x"58",
          4419 => x"80",
          4420 => x"06",
          4421 => x"06",
          4422 => x"19",
          4423 => x"57",
          4424 => x"b9",
          4425 => x"b6",
          4426 => x"e0",
          4427 => x"84",
          4428 => x"33",
          4429 => x"05",
          4430 => x"70",
          4431 => x"33",
          4432 => x"05",
          4433 => x"15",
          4434 => x"33",
          4435 => x"33",
          4436 => x"19",
          4437 => x"55",
          4438 => x"ce",
          4439 => x"72",
          4440 => x"0c",
          4441 => x"04",
          4442 => x"94",
          4443 => x"92",
          4444 => x"ff",
          4445 => x"b6",
          4446 => x"55",
          4447 => x"27",
          4448 => x"77",
          4449 => x"dd",
          4450 => x"ff",
          4451 => x"83",
          4452 => x"56",
          4453 => x"2e",
          4454 => x"fe",
          4455 => x"76",
          4456 => x"84",
          4457 => x"71",
          4458 => x"72",
          4459 => x"52",
          4460 => x"73",
          4461 => x"38",
          4462 => x"33",
          4463 => x"15",
          4464 => x"55",
          4465 => x"0b",
          4466 => x"34",
          4467 => x"81",
          4468 => x"ff",
          4469 => x"80",
          4470 => x"38",
          4471 => x"e0",
          4472 => x"75",
          4473 => x"57",
          4474 => x"53",
          4475 => x"fd",
          4476 => x"0b",
          4477 => x"33",
          4478 => x"89",
          4479 => x"96",
          4480 => x"84",
          4481 => x"33",
          4482 => x"b6",
          4483 => x"fc",
          4484 => x"3d",
          4485 => x"84",
          4486 => x"33",
          4487 => x"86",
          4488 => x"70",
          4489 => x"c3",
          4490 => x"70",
          4491 => x"b6",
          4492 => x"71",
          4493 => x"38",
          4494 => x"95",
          4495 => x"84",
          4496 => x"86",
          4497 => x"80",
          4498 => x"95",
          4499 => x"94",
          4500 => x"ff",
          4501 => x"72",
          4502 => x"38",
          4503 => x"70",
          4504 => x"34",
          4505 => x"b8",
          4506 => x"3d",
          4507 => x"f8",
          4508 => x"73",
          4509 => x"70",
          4510 => x"06",
          4511 => x"54",
          4512 => x"94",
          4513 => x"83",
          4514 => x"72",
          4515 => x"d7",
          4516 => x"55",
          4517 => x"75",
          4518 => x"70",
          4519 => x"f8",
          4520 => x"0b",
          4521 => x"0c",
          4522 => x"04",
          4523 => x"33",
          4524 => x"70",
          4525 => x"2c",
          4526 => x"56",
          4527 => x"83",
          4528 => x"80",
          4529 => x"e4",
          4530 => x"0d",
          4531 => x"95",
          4532 => x"84",
          4533 => x"ff",
          4534 => x"51",
          4535 => x"83",
          4536 => x"72",
          4537 => x"34",
          4538 => x"b8",
          4539 => x"3d",
          4540 => x"0b",
          4541 => x"34",
          4542 => x"33",
          4543 => x"33",
          4544 => x"52",
          4545 => x"fe",
          4546 => x"12",
          4547 => x"f8",
          4548 => x"d0",
          4549 => x"0d",
          4550 => x"33",
          4551 => x"26",
          4552 => x"10",
          4553 => x"f8",
          4554 => x"08",
          4555 => x"90",
          4556 => x"f0",
          4557 => x"2b",
          4558 => x"70",
          4559 => x"07",
          4560 => x"51",
          4561 => x"2e",
          4562 => x"9c",
          4563 => x"0b",
          4564 => x"34",
          4565 => x"b8",
          4566 => x"3d",
          4567 => x"f8",
          4568 => x"9f",
          4569 => x"51",
          4570 => x"90",
          4571 => x"84",
          4572 => x"83",
          4573 => x"83",
          4574 => x"80",
          4575 => x"70",
          4576 => x"34",
          4577 => x"f8",
          4578 => x"fe",
          4579 => x"51",
          4580 => x"90",
          4581 => x"80",
          4582 => x"f8",
          4583 => x"0b",
          4584 => x"0c",
          4585 => x"04",
          4586 => x"33",
          4587 => x"84",
          4588 => x"83",
          4589 => x"ff",
          4590 => x"f8",
          4591 => x"07",
          4592 => x"f8",
          4593 => x"a5",
          4594 => x"90",
          4595 => x"06",
          4596 => x"70",
          4597 => x"34",
          4598 => x"83",
          4599 => x"81",
          4600 => x"07",
          4601 => x"f8",
          4602 => x"81",
          4603 => x"90",
          4604 => x"06",
          4605 => x"70",
          4606 => x"34",
          4607 => x"83",
          4608 => x"81",
          4609 => x"70",
          4610 => x"34",
          4611 => x"83",
          4612 => x"81",
          4613 => x"d0",
          4614 => x"83",
          4615 => x"fe",
          4616 => x"f8",
          4617 => x"bf",
          4618 => x"51",
          4619 => x"90",
          4620 => x"39",
          4621 => x"33",
          4622 => x"80",
          4623 => x"70",
          4624 => x"34",
          4625 => x"83",
          4626 => x"81",
          4627 => x"c0",
          4628 => x"83",
          4629 => x"fe",
          4630 => x"f8",
          4631 => x"af",
          4632 => x"51",
          4633 => x"90",
          4634 => x"39",
          4635 => x"33",
          4636 => x"51",
          4637 => x"90",
          4638 => x"39",
          4639 => x"33",
          4640 => x"82",
          4641 => x"83",
          4642 => x"fd",
          4643 => x"3d",
          4644 => x"05",
          4645 => x"05",
          4646 => x"33",
          4647 => x"33",
          4648 => x"33",
          4649 => x"33",
          4650 => x"33",
          4651 => x"5d",
          4652 => x"82",
          4653 => x"38",
          4654 => x"a5",
          4655 => x"2e",
          4656 => x"7d",
          4657 => x"34",
          4658 => x"b6",
          4659 => x"83",
          4660 => x"7b",
          4661 => x"23",
          4662 => x"95",
          4663 => x"0d",
          4664 => x"2e",
          4665 => x"db",
          4666 => x"84",
          4667 => x"81",
          4668 => x"dc",
          4669 => x"83",
          4670 => x"a8",
          4671 => x"95",
          4672 => x"83",
          4673 => x"79",
          4674 => x"d8",
          4675 => x"b6",
          4676 => x"84",
          4677 => x"55",
          4678 => x"53",
          4679 => x"e2",
          4680 => x"81",
          4681 => x"84",
          4682 => x"80",
          4683 => x"dc",
          4684 => x"f8",
          4685 => x"83",
          4686 => x"7c",
          4687 => x"34",
          4688 => x"04",
          4689 => x"b6",
          4690 => x"0b",
          4691 => x"34",
          4692 => x"f8",
          4693 => x"0b",
          4694 => x"34",
          4695 => x"f8",
          4696 => x"b7",
          4697 => x"84",
          4698 => x"57",
          4699 => x"33",
          4700 => x"7b",
          4701 => x"7a",
          4702 => x"f4",
          4703 => x"8b",
          4704 => x"84",
          4705 => x"5a",
          4706 => x"27",
          4707 => x"10",
          4708 => x"05",
          4709 => x"59",
          4710 => x"51",
          4711 => x"3f",
          4712 => x"81",
          4713 => x"b7",
          4714 => x"5b",
          4715 => x"26",
          4716 => x"d2",
          4717 => x"80",
          4718 => x"84",
          4719 => x"80",
          4720 => x"dc",
          4721 => x"f8",
          4722 => x"83",
          4723 => x"7c",
          4724 => x"34",
          4725 => x"04",
          4726 => x"b6",
          4727 => x"0b",
          4728 => x"34",
          4729 => x"f8",
          4730 => x"0b",
          4731 => x"34",
          4732 => x"f8",
          4733 => x"f6",
          4734 => x"92",
          4735 => x"b8",
          4736 => x"83",
          4737 => x"ff",
          4738 => x"80",
          4739 => x"c8",
          4740 => x"97",
          4741 => x"b8",
          4742 => x"fd",
          4743 => x"f6",
          4744 => x"52",
          4745 => x"51",
          4746 => x"3f",
          4747 => x"81",
          4748 => x"5a",
          4749 => x"3d",
          4750 => x"84",
          4751 => x"33",
          4752 => x"33",
          4753 => x"33",
          4754 => x"33",
          4755 => x"12",
          4756 => x"80",
          4757 => x"92",
          4758 => x"59",
          4759 => x"29",
          4760 => x"ff",
          4761 => x"f6",
          4762 => x"59",
          4763 => x"57",
          4764 => x"81",
          4765 => x"89",
          4766 => x"38",
          4767 => x"81",
          4768 => x"81",
          4769 => x"38",
          4770 => x"82",
          4771 => x"b6",
          4772 => x"f8",
          4773 => x"f8",
          4774 => x"72",
          4775 => x"56",
          4776 => x"e0",
          4777 => x"a7",
          4778 => x"34",
          4779 => x"33",
          4780 => x"33",
          4781 => x"22",
          4782 => x"12",
          4783 => x"53",
          4784 => x"96",
          4785 => x"f8",
          4786 => x"71",
          4787 => x"54",
          4788 => x"33",
          4789 => x"80",
          4790 => x"b6",
          4791 => x"81",
          4792 => x"f8",
          4793 => x"f8",
          4794 => x"72",
          4795 => x"5b",
          4796 => x"83",
          4797 => x"84",
          4798 => x"34",
          4799 => x"81",
          4800 => x"55",
          4801 => x"81",
          4802 => x"b6",
          4803 => x"77",
          4804 => x"ff",
          4805 => x"83",
          4806 => x"84",
          4807 => x"53",
          4808 => x"8c",
          4809 => x"dc",
          4810 => x"80",
          4811 => x"38",
          4812 => x"b8",
          4813 => x"3d",
          4814 => x"8d",
          4815 => x"75",
          4816 => x"f7",
          4817 => x"2e",
          4818 => x"fe",
          4819 => x"52",
          4820 => x"96",
          4821 => x"83",
          4822 => x"ff",
          4823 => x"f8",
          4824 => x"53",
          4825 => x"13",
          4826 => x"75",
          4827 => x"81",
          4828 => x"38",
          4829 => x"52",
          4830 => x"ba",
          4831 => x"70",
          4832 => x"54",
          4833 => x"26",
          4834 => x"76",
          4835 => x"fd",
          4836 => x"13",
          4837 => x"06",
          4838 => x"73",
          4839 => x"fe",
          4840 => x"83",
          4841 => x"fe",
          4842 => x"52",
          4843 => x"de",
          4844 => x"84",
          4845 => x"89",
          4846 => x"75",
          4847 => x"09",
          4848 => x"ca",
          4849 => x"95",
          4850 => x"ff",
          4851 => x"05",
          4852 => x"38",
          4853 => x"83",
          4854 => x"76",
          4855 => x"fc",
          4856 => x"f8",
          4857 => x"81",
          4858 => x"ff",
          4859 => x"fe",
          4860 => x"53",
          4861 => x"95",
          4862 => x"39",
          4863 => x"f8",
          4864 => x"52",
          4865 => x"e2",
          4866 => x"39",
          4867 => x"51",
          4868 => x"fe",
          4869 => x"3d",
          4870 => x"f3",
          4871 => x"b7",
          4872 => x"59",
          4873 => x"81",
          4874 => x"82",
          4875 => x"38",
          4876 => x"84",
          4877 => x"8a",
          4878 => x"38",
          4879 => x"84",
          4880 => x"89",
          4881 => x"38",
          4882 => x"33",
          4883 => x"33",
          4884 => x"33",
          4885 => x"05",
          4886 => x"84",
          4887 => x"33",
          4888 => x"80",
          4889 => x"b6",
          4890 => x"f8",
          4891 => x"f8",
          4892 => x"71",
          4893 => x"5a",
          4894 => x"83",
          4895 => x"34",
          4896 => x"33",
          4897 => x"62",
          4898 => x"83",
          4899 => x"7f",
          4900 => x"80",
          4901 => x"b6",
          4902 => x"81",
          4903 => x"f8",
          4904 => x"f8",
          4905 => x"72",
          4906 => x"40",
          4907 => x"83",
          4908 => x"84",
          4909 => x"34",
          4910 => x"81",
          4911 => x"58",
          4912 => x"81",
          4913 => x"b6",
          4914 => x"79",
          4915 => x"ff",
          4916 => x"83",
          4917 => x"80",
          4918 => x"e4",
          4919 => x"0d",
          4920 => x"2e",
          4921 => x"b7",
          4922 => x"fd",
          4923 => x"2e",
          4924 => x"78",
          4925 => x"89",
          4926 => x"0b",
          4927 => x"0c",
          4928 => x"33",
          4929 => x"33",
          4930 => x"33",
          4931 => x"05",
          4932 => x"84",
          4933 => x"33",
          4934 => x"80",
          4935 => x"b6",
          4936 => x"f8",
          4937 => x"f8",
          4938 => x"71",
          4939 => x"5f",
          4940 => x"83",
          4941 => x"34",
          4942 => x"33",
          4943 => x"19",
          4944 => x"f8",
          4945 => x"a7",
          4946 => x"34",
          4947 => x"33",
          4948 => x"06",
          4949 => x"22",
          4950 => x"33",
          4951 => x"11",
          4952 => x"58",
          4953 => x"90",
          4954 => x"97",
          4955 => x"81",
          4956 => x"81",
          4957 => x"60",
          4958 => x"ca",
          4959 => x"f8",
          4960 => x"0b",
          4961 => x"0c",
          4962 => x"04",
          4963 => x"82",
          4964 => x"9b",
          4965 => x"38",
          4966 => x"09",
          4967 => x"a8",
          4968 => x"83",
          4969 => x"80",
          4970 => x"e4",
          4971 => x"0d",
          4972 => x"2e",
          4973 => x"d0",
          4974 => x"89",
          4975 => x"38",
          4976 => x"33",
          4977 => x"57",
          4978 => x"e4",
          4979 => x"b7",
          4980 => x"77",
          4981 => x"59",
          4982 => x"b7",
          4983 => x"80",
          4984 => x"e4",
          4985 => x"0d",
          4986 => x"2e",
          4987 => x"80",
          4988 => x"e0",
          4989 => x"d8",
          4990 => x"94",
          4991 => x"95",
          4992 => x"29",
          4993 => x"40",
          4994 => x"19",
          4995 => x"a0",
          4996 => x"84",
          4997 => x"83",
          4998 => x"83",
          4999 => x"72",
          5000 => x"41",
          5001 => x"78",
          5002 => x"1f",
          5003 => x"94",
          5004 => x"29",
          5005 => x"83",
          5006 => x"86",
          5007 => x"1b",
          5008 => x"d8",
          5009 => x"ff",
          5010 => x"92",
          5011 => x"95",
          5012 => x"29",
          5013 => x"43",
          5014 => x"f8",
          5015 => x"84",
          5016 => x"34",
          5017 => x"fe",
          5018 => x"52",
          5019 => x"fa",
          5020 => x"83",
          5021 => x"fe",
          5022 => x"b6",
          5023 => x"f8",
          5024 => x"81",
          5025 => x"f8",
          5026 => x"71",
          5027 => x"a7",
          5028 => x"83",
          5029 => x"40",
          5030 => x"7e",
          5031 => x"83",
          5032 => x"83",
          5033 => x"5a",
          5034 => x"5c",
          5035 => x"86",
          5036 => x"81",
          5037 => x"1a",
          5038 => x"fc",
          5039 => x"56",
          5040 => x"95",
          5041 => x"39",
          5042 => x"b7",
          5043 => x"0b",
          5044 => x"34",
          5045 => x"b7",
          5046 => x"0b",
          5047 => x"34",
          5048 => x"b7",
          5049 => x"0b",
          5050 => x"0c",
          5051 => x"04",
          5052 => x"33",
          5053 => x"34",
          5054 => x"33",
          5055 => x"34",
          5056 => x"33",
          5057 => x"34",
          5058 => x"b7",
          5059 => x"0b",
          5060 => x"0c",
          5061 => x"04",
          5062 => x"2e",
          5063 => x"fa",
          5064 => x"f8",
          5065 => x"b6",
          5066 => x"81",
          5067 => x"f8",
          5068 => x"81",
          5069 => x"75",
          5070 => x"a7",
          5071 => x"83",
          5072 => x"5c",
          5073 => x"29",
          5074 => x"ff",
          5075 => x"f6",
          5076 => x"5c",
          5077 => x"5b",
          5078 => x"2e",
          5079 => x"78",
          5080 => x"ff",
          5081 => x"75",
          5082 => x"57",
          5083 => x"95",
          5084 => x"ff",
          5085 => x"ff",
          5086 => x"ff",
          5087 => x"29",
          5088 => x"5b",
          5089 => x"33",
          5090 => x"80",
          5091 => x"b6",
          5092 => x"f8",
          5093 => x"f8",
          5094 => x"71",
          5095 => x"5e",
          5096 => x"0b",
          5097 => x"18",
          5098 => x"94",
          5099 => x"29",
          5100 => x"56",
          5101 => x"33",
          5102 => x"80",
          5103 => x"b6",
          5104 => x"81",
          5105 => x"f8",
          5106 => x"f8",
          5107 => x"72",
          5108 => x"5d",
          5109 => x"83",
          5110 => x"7f",
          5111 => x"05",
          5112 => x"70",
          5113 => x"5c",
          5114 => x"26",
          5115 => x"84",
          5116 => x"5a",
          5117 => x"38",
          5118 => x"77",
          5119 => x"34",
          5120 => x"33",
          5121 => x"06",
          5122 => x"56",
          5123 => x"78",
          5124 => x"d8",
          5125 => x"2e",
          5126 => x"78",
          5127 => x"a8",
          5128 => x"e4",
          5129 => x"83",
          5130 => x"bf",
          5131 => x"b4",
          5132 => x"38",
          5133 => x"83",
          5134 => x"58",
          5135 => x"80",
          5136 => x"95",
          5137 => x"81",
          5138 => x"3f",
          5139 => x"b8",
          5140 => x"3d",
          5141 => x"f8",
          5142 => x"b6",
          5143 => x"81",
          5144 => x"f8",
          5145 => x"81",
          5146 => x"75",
          5147 => x"a7",
          5148 => x"83",
          5149 => x"5c",
          5150 => x"29",
          5151 => x"ff",
          5152 => x"f6",
          5153 => x"53",
          5154 => x"5b",
          5155 => x"2e",
          5156 => x"80",
          5157 => x"ff",
          5158 => x"ff",
          5159 => x"ff",
          5160 => x"29",
          5161 => x"40",
          5162 => x"33",
          5163 => x"80",
          5164 => x"b6",
          5165 => x"f8",
          5166 => x"f8",
          5167 => x"71",
          5168 => x"41",
          5169 => x"0b",
          5170 => x"1c",
          5171 => x"94",
          5172 => x"29",
          5173 => x"83",
          5174 => x"86",
          5175 => x"1a",
          5176 => x"d8",
          5177 => x"ff",
          5178 => x"92",
          5179 => x"95",
          5180 => x"29",
          5181 => x"5a",
          5182 => x"f8",
          5183 => x"97",
          5184 => x"60",
          5185 => x"81",
          5186 => x"58",
          5187 => x"81",
          5188 => x"b6",
          5189 => x"77",
          5190 => x"ff",
          5191 => x"83",
          5192 => x"81",
          5193 => x"ff",
          5194 => x"7b",
          5195 => x"a7",
          5196 => x"94",
          5197 => x"d8",
          5198 => x"95",
          5199 => x"ff",
          5200 => x"ff",
          5201 => x"ff",
          5202 => x"29",
          5203 => x"43",
          5204 => x"84",
          5205 => x"86",
          5206 => x"1b",
          5207 => x"d8",
          5208 => x"95",
          5209 => x"92",
          5210 => x"29",
          5211 => x"5e",
          5212 => x"83",
          5213 => x"34",
          5214 => x"33",
          5215 => x"1e",
          5216 => x"f8",
          5217 => x"a7",
          5218 => x"34",
          5219 => x"33",
          5220 => x"06",
          5221 => x"22",
          5222 => x"33",
          5223 => x"11",
          5224 => x"40",
          5225 => x"90",
          5226 => x"b6",
          5227 => x"81",
          5228 => x"ff",
          5229 => x"79",
          5230 => x"d6",
          5231 => x"f8",
          5232 => x"df",
          5233 => x"84",
          5234 => x"80",
          5235 => x"e4",
          5236 => x"0d",
          5237 => x"96",
          5238 => x"84",
          5239 => x"33",
          5240 => x"f8",
          5241 => x"81",
          5242 => x"ff",
          5243 => x"ca",
          5244 => x"84",
          5245 => x"80",
          5246 => x"e4",
          5247 => x"0d",
          5248 => x"96",
          5249 => x"84",
          5250 => x"33",
          5251 => x"f8",
          5252 => x"b6",
          5253 => x"f8",
          5254 => x"5b",
          5255 => x"fc",
          5256 => x"b7",
          5257 => x"3d",
          5258 => x"d8",
          5259 => x"8a",
          5260 => x"b8",
          5261 => x"2e",
          5262 => x"84",
          5263 => x"81",
          5264 => x"75",
          5265 => x"34",
          5266 => x"fe",
          5267 => x"80",
          5268 => x"61",
          5269 => x"05",
          5270 => x"39",
          5271 => x"17",
          5272 => x"b6",
          5273 => x"7b",
          5274 => x"94",
          5275 => x"d8",
          5276 => x"95",
          5277 => x"5c",
          5278 => x"84",
          5279 => x"83",
          5280 => x"83",
          5281 => x"72",
          5282 => x"41",
          5283 => x"b6",
          5284 => x"7f",
          5285 => x"80",
          5286 => x"b6",
          5287 => x"f8",
          5288 => x"f8",
          5289 => x"71",
          5290 => x"43",
          5291 => x"83",
          5292 => x"34",
          5293 => x"33",
          5294 => x"1b",
          5295 => x"f8",
          5296 => x"86",
          5297 => x"05",
          5298 => x"d8",
          5299 => x"ff",
          5300 => x"92",
          5301 => x"95",
          5302 => x"29",
          5303 => x"5a",
          5304 => x"f8",
          5305 => x"97",
          5306 => x"81",
          5307 => x"ff",
          5308 => x"60",
          5309 => x"a2",
          5310 => x"d9",
          5311 => x"90",
          5312 => x"1a",
          5313 => x"f8",
          5314 => x"0b",
          5315 => x"0c",
          5316 => x"33",
          5317 => x"2e",
          5318 => x"84",
          5319 => x"56",
          5320 => x"38",
          5321 => x"51",
          5322 => x"80",
          5323 => x"e4",
          5324 => x"0d",
          5325 => x"cc",
          5326 => x"94",
          5327 => x"cd",
          5328 => x"95",
          5329 => x"ce",
          5330 => x"83",
          5331 => x"ff",
          5332 => x"f8",
          5333 => x"b8",
          5334 => x"f8",
          5335 => x"b8",
          5336 => x"f8",
          5337 => x"b8",
          5338 => x"9e",
          5339 => x"e5",
          5340 => x"80",
          5341 => x"38",
          5342 => x"22",
          5343 => x"2e",
          5344 => x"ff",
          5345 => x"f8",
          5346 => x"05",
          5347 => x"94",
          5348 => x"54",
          5349 => x"e3",
          5350 => x"3d",
          5351 => x"fe",
          5352 => x"76",
          5353 => x"83",
          5354 => x"e4",
          5355 => x"06",
          5356 => x"33",
          5357 => x"41",
          5358 => x"fe",
          5359 => x"52",
          5360 => x"51",
          5361 => x"3f",
          5362 => x"80",
          5363 => x"e5",
          5364 => x"79",
          5365 => x"5b",
          5366 => x"fe",
          5367 => x"10",
          5368 => x"05",
          5369 => x"57",
          5370 => x"26",
          5371 => x"75",
          5372 => x"c7",
          5373 => x"7e",
          5374 => x"b7",
          5375 => x"7d",
          5376 => x"a4",
          5377 => x"94",
          5378 => x"b9",
          5379 => x"31",
          5380 => x"9f",
          5381 => x"5a",
          5382 => x"5c",
          5383 => x"94",
          5384 => x"39",
          5385 => x"33",
          5386 => x"2e",
          5387 => x"84",
          5388 => x"ff",
          5389 => x"ff",
          5390 => x"d8",
          5391 => x"5f",
          5392 => x"fd",
          5393 => x"83",
          5394 => x"fd",
          5395 => x"0b",
          5396 => x"34",
          5397 => x"33",
          5398 => x"06",
          5399 => x"80",
          5400 => x"38",
          5401 => x"75",
          5402 => x"34",
          5403 => x"80",
          5404 => x"95",
          5405 => x"94",
          5406 => x"d7",
          5407 => x"57",
          5408 => x"25",
          5409 => x"81",
          5410 => x"83",
          5411 => x"fc",
          5412 => x"b7",
          5413 => x"7f",
          5414 => x"e0",
          5415 => x"95",
          5416 => x"b9",
          5417 => x"31",
          5418 => x"9f",
          5419 => x"5a",
          5420 => x"5a",
          5421 => x"95",
          5422 => x"39",
          5423 => x"33",
          5424 => x"2e",
          5425 => x"84",
          5426 => x"41",
          5427 => x"09",
          5428 => x"b6",
          5429 => x"d8",
          5430 => x"95",
          5431 => x"94",
          5432 => x"29",
          5433 => x"a0",
          5434 => x"f8",
          5435 => x"51",
          5436 => x"60",
          5437 => x"83",
          5438 => x"83",
          5439 => x"87",
          5440 => x"06",
          5441 => x"5d",
          5442 => x"80",
          5443 => x"38",
          5444 => x"f6",
          5445 => x"f2",
          5446 => x"e5",
          5447 => x"80",
          5448 => x"38",
          5449 => x"22",
          5450 => x"2e",
          5451 => x"fb",
          5452 => x"0b",
          5453 => x"34",
          5454 => x"84",
          5455 => x"56",
          5456 => x"90",
          5457 => x"b8",
          5458 => x"f8",
          5459 => x"7c",
          5460 => x"d8",
          5461 => x"59",
          5462 => x"7d",
          5463 => x"75",
          5464 => x"f8",
          5465 => x"a2",
          5466 => x"e5",
          5467 => x"80",
          5468 => x"38",
          5469 => x"33",
          5470 => x"33",
          5471 => x"84",
          5472 => x"ff",
          5473 => x"56",
          5474 => x"83",
          5475 => x"76",
          5476 => x"34",
          5477 => x"83",
          5478 => x"fe",
          5479 => x"80",
          5480 => x"e5",
          5481 => x"76",
          5482 => x"c7",
          5483 => x"84",
          5484 => x"70",
          5485 => x"83",
          5486 => x"fe",
          5487 => x"81",
          5488 => x"ff",
          5489 => x"e5",
          5490 => x"58",
          5491 => x"0b",
          5492 => x"33",
          5493 => x"80",
          5494 => x"84",
          5495 => x"56",
          5496 => x"83",
          5497 => x"81",
          5498 => x"ff",
          5499 => x"f3",
          5500 => x"39",
          5501 => x"33",
          5502 => x"27",
          5503 => x"84",
          5504 => x"ff",
          5505 => x"ff",
          5506 => x"b9",
          5507 => x"70",
          5508 => x"84",
          5509 => x"70",
          5510 => x"ff",
          5511 => x"52",
          5512 => x"5c",
          5513 => x"83",
          5514 => x"79",
          5515 => x"23",
          5516 => x"06",
          5517 => x"5f",
          5518 => x"83",
          5519 => x"76",
          5520 => x"34",
          5521 => x"33",
          5522 => x"40",
          5523 => x"f9",
          5524 => x"56",
          5525 => x"95",
          5526 => x"39",
          5527 => x"33",
          5528 => x"2e",
          5529 => x"84",
          5530 => x"84",
          5531 => x"40",
          5532 => x"26",
          5533 => x"83",
          5534 => x"84",
          5535 => x"70",
          5536 => x"83",
          5537 => x"71",
          5538 => x"86",
          5539 => x"05",
          5540 => x"22",
          5541 => x"7e",
          5542 => x"83",
          5543 => x"83",
          5544 => x"46",
          5545 => x"5f",
          5546 => x"2e",
          5547 => x"79",
          5548 => x"06",
          5549 => x"5d",
          5550 => x"24",
          5551 => x"84",
          5552 => x"56",
          5553 => x"8e",
          5554 => x"16",
          5555 => x"f8",
          5556 => x"81",
          5557 => x"7c",
          5558 => x"80",
          5559 => x"e5",
          5560 => x"d7",
          5561 => x"76",
          5562 => x"38",
          5563 => x"75",
          5564 => x"34",
          5565 => x"06",
          5566 => x"22",
          5567 => x"5a",
          5568 => x"90",
          5569 => x"31",
          5570 => x"81",
          5571 => x"71",
          5572 => x"5b",
          5573 => x"a7",
          5574 => x"86",
          5575 => x"7f",
          5576 => x"7f",
          5577 => x"71",
          5578 => x"42",
          5579 => x"79",
          5580 => x"d6",
          5581 => x"b6",
          5582 => x"e0",
          5583 => x"84",
          5584 => x"33",
          5585 => x"05",
          5586 => x"70",
          5587 => x"33",
          5588 => x"05",
          5589 => x"18",
          5590 => x"33",
          5591 => x"33",
          5592 => x"1d",
          5593 => x"58",
          5594 => x"f7",
          5595 => x"e0",
          5596 => x"84",
          5597 => x"33",
          5598 => x"05",
          5599 => x"70",
          5600 => x"33",
          5601 => x"05",
          5602 => x"18",
          5603 => x"33",
          5604 => x"33",
          5605 => x"1d",
          5606 => x"58",
          5607 => x"ff",
          5608 => x"e6",
          5609 => x"e5",
          5610 => x"80",
          5611 => x"38",
          5612 => x"b8",
          5613 => x"d8",
          5614 => x"ce",
          5615 => x"84",
          5616 => x"ff",
          5617 => x"e5",
          5618 => x"40",
          5619 => x"2e",
          5620 => x"b8",
          5621 => x"75",
          5622 => x"81",
          5623 => x"38",
          5624 => x"33",
          5625 => x"ff",
          5626 => x"94",
          5627 => x"5c",
          5628 => x"2e",
          5629 => x"84",
          5630 => x"40",
          5631 => x"f6",
          5632 => x"81",
          5633 => x"60",
          5634 => x"fe",
          5635 => x"26",
          5636 => x"07",
          5637 => x"f2",
          5638 => x"10",
          5639 => x"29",
          5640 => x"a7",
          5641 => x"70",
          5642 => x"86",
          5643 => x"05",
          5644 => x"58",
          5645 => x"8b",
          5646 => x"83",
          5647 => x"8b",
          5648 => x"f8",
          5649 => x"98",
          5650 => x"2b",
          5651 => x"2b",
          5652 => x"79",
          5653 => x"5f",
          5654 => x"27",
          5655 => x"77",
          5656 => x"59",
          5657 => x"70",
          5658 => x"0c",
          5659 => x"ee",
          5660 => x"d8",
          5661 => x"d7",
          5662 => x"7e",
          5663 => x"60",
          5664 => x"83",
          5665 => x"7d",
          5666 => x"05",
          5667 => x"5a",
          5668 => x"8c",
          5669 => x"31",
          5670 => x"29",
          5671 => x"40",
          5672 => x"57",
          5673 => x"26",
          5674 => x"83",
          5675 => x"84",
          5676 => x"59",
          5677 => x"e0",
          5678 => x"79",
          5679 => x"05",
          5680 => x"17",
          5681 => x"26",
          5682 => x"a0",
          5683 => x"19",
          5684 => x"70",
          5685 => x"34",
          5686 => x"75",
          5687 => x"38",
          5688 => x"ff",
          5689 => x"ff",
          5690 => x"fe",
          5691 => x"f8",
          5692 => x"80",
          5693 => x"84",
          5694 => x"06",
          5695 => x"07",
          5696 => x"7b",
          5697 => x"09",
          5698 => x"38",
          5699 => x"83",
          5700 => x"81",
          5701 => x"ff",
          5702 => x"f5",
          5703 => x"f8",
          5704 => x"5e",
          5705 => x"1e",
          5706 => x"83",
          5707 => x"84",
          5708 => x"83",
          5709 => x"84",
          5710 => x"42",
          5711 => x"fa",
          5712 => x"f8",
          5713 => x"07",
          5714 => x"f8",
          5715 => x"18",
          5716 => x"06",
          5717 => x"fb",
          5718 => x"90",
          5719 => x"06",
          5720 => x"75",
          5721 => x"34",
          5722 => x"f8",
          5723 => x"fb",
          5724 => x"56",
          5725 => x"90",
          5726 => x"83",
          5727 => x"81",
          5728 => x"07",
          5729 => x"f8",
          5730 => x"39",
          5731 => x"33",
          5732 => x"90",
          5733 => x"83",
          5734 => x"ff",
          5735 => x"f1",
          5736 => x"90",
          5737 => x"70",
          5738 => x"59",
          5739 => x"39",
          5740 => x"33",
          5741 => x"56",
          5742 => x"90",
          5743 => x"39",
          5744 => x"33",
          5745 => x"90",
          5746 => x"83",
          5747 => x"fe",
          5748 => x"f8",
          5749 => x"ef",
          5750 => x"07",
          5751 => x"f8",
          5752 => x"ea",
          5753 => x"90",
          5754 => x"06",
          5755 => x"56",
          5756 => x"90",
          5757 => x"39",
          5758 => x"33",
          5759 => x"a0",
          5760 => x"83",
          5761 => x"fe",
          5762 => x"f8",
          5763 => x"fe",
          5764 => x"56",
          5765 => x"90",
          5766 => x"39",
          5767 => x"33",
          5768 => x"84",
          5769 => x"83",
          5770 => x"fe",
          5771 => x"f8",
          5772 => x"fa",
          5773 => x"56",
          5774 => x"90",
          5775 => x"39",
          5776 => x"33",
          5777 => x"56",
          5778 => x"90",
          5779 => x"39",
          5780 => x"33",
          5781 => x"56",
          5782 => x"90",
          5783 => x"39",
          5784 => x"33",
          5785 => x"56",
          5786 => x"90",
          5787 => x"39",
          5788 => x"33",
          5789 => x"80",
          5790 => x"75",
          5791 => x"34",
          5792 => x"83",
          5793 => x"81",
          5794 => x"07",
          5795 => x"f8",
          5796 => x"ba",
          5797 => x"83",
          5798 => x"80",
          5799 => x"d2",
          5800 => x"ff",
          5801 => x"cc",
          5802 => x"94",
          5803 => x"cd",
          5804 => x"95",
          5805 => x"ce",
          5806 => x"83",
          5807 => x"80",
          5808 => x"e0",
          5809 => x"39",
          5810 => x"b7",
          5811 => x"0b",
          5812 => x"0c",
          5813 => x"04",
          5814 => x"95",
          5815 => x"95",
          5816 => x"ff",
          5817 => x"05",
          5818 => x"39",
          5819 => x"42",
          5820 => x"11",
          5821 => x"51",
          5822 => x"3f",
          5823 => x"08",
          5824 => x"b8",
          5825 => x"b7",
          5826 => x"0b",
          5827 => x"34",
          5828 => x"b8",
          5829 => x"3d",
          5830 => x"83",
          5831 => x"ef",
          5832 => x"b7",
          5833 => x"11",
          5834 => x"84",
          5835 => x"7b",
          5836 => x"06",
          5837 => x"ca",
          5838 => x"b8",
          5839 => x"80",
          5840 => x"e4",
          5841 => x"80",
          5842 => x"95",
          5843 => x"81",
          5844 => x"3f",
          5845 => x"33",
          5846 => x"06",
          5847 => x"56",
          5848 => x"80",
          5849 => x"95",
          5850 => x"81",
          5851 => x"3f",
          5852 => x"8a",
          5853 => x"e9",
          5854 => x"39",
          5855 => x"33",
          5856 => x"09",
          5857 => x"72",
          5858 => x"57",
          5859 => x"75",
          5860 => x"d9",
          5861 => x"d8",
          5862 => x"60",
          5863 => x"38",
          5864 => x"95",
          5865 => x"39",
          5866 => x"33",
          5867 => x"09",
          5868 => x"72",
          5869 => x"57",
          5870 => x"83",
          5871 => x"81",
          5872 => x"d7",
          5873 => x"59",
          5874 => x"78",
          5875 => x"38",
          5876 => x"bb",
          5877 => x"d7",
          5878 => x"ff",
          5879 => x"81",
          5880 => x"a6",
          5881 => x"94",
          5882 => x"d8",
          5883 => x"ff",
          5884 => x"95",
          5885 => x"29",
          5886 => x"a0",
          5887 => x"f8",
          5888 => x"5f",
          5889 => x"05",
          5890 => x"ff",
          5891 => x"ea",
          5892 => x"44",
          5893 => x"77",
          5894 => x"f5",
          5895 => x"ff",
          5896 => x"11",
          5897 => x"7b",
          5898 => x"38",
          5899 => x"33",
          5900 => x"27",
          5901 => x"ff",
          5902 => x"83",
          5903 => x"7c",
          5904 => x"ff",
          5905 => x"80",
          5906 => x"df",
          5907 => x"d7",
          5908 => x"76",
          5909 => x"38",
          5910 => x"75",
          5911 => x"34",
          5912 => x"06",
          5913 => x"22",
          5914 => x"5a",
          5915 => x"90",
          5916 => x"31",
          5917 => x"81",
          5918 => x"71",
          5919 => x"5f",
          5920 => x"a7",
          5921 => x"86",
          5922 => x"7c",
          5923 => x"7f",
          5924 => x"71",
          5925 => x"41",
          5926 => x"79",
          5927 => x"ea",
          5928 => x"b6",
          5929 => x"e0",
          5930 => x"84",
          5931 => x"33",
          5932 => x"05",
          5933 => x"70",
          5934 => x"33",
          5935 => x"05",
          5936 => x"18",
          5937 => x"33",
          5938 => x"33",
          5939 => x"1d",
          5940 => x"58",
          5941 => x"ec",
          5942 => x"e0",
          5943 => x"84",
          5944 => x"33",
          5945 => x"05",
          5946 => x"70",
          5947 => x"33",
          5948 => x"05",
          5949 => x"18",
          5950 => x"33",
          5951 => x"33",
          5952 => x"1d",
          5953 => x"58",
          5954 => x"ff",
          5955 => x"fa",
          5956 => x"96",
          5957 => x"84",
          5958 => x"33",
          5959 => x"f8",
          5960 => x"b6",
          5961 => x"f8",
          5962 => x"b6",
          5963 => x"5c",
          5964 => x"e9",
          5965 => x"d2",
          5966 => x"d7",
          5967 => x"ff",
          5968 => x"5c",
          5969 => x"61",
          5970 => x"76",
          5971 => x"f8",
          5972 => x"81",
          5973 => x"19",
          5974 => x"7a",
          5975 => x"80",
          5976 => x"f8",
          5977 => x"b6",
          5978 => x"81",
          5979 => x"12",
          5980 => x"80",
          5981 => x"8d",
          5982 => x"75",
          5983 => x"34",
          5984 => x"83",
          5985 => x"81",
          5986 => x"d8",
          5987 => x"59",
          5988 => x"7f",
          5989 => x"38",
          5990 => x"c5",
          5991 => x"2e",
          5992 => x"f4",
          5993 => x"f8",
          5994 => x"81",
          5995 => x"f8",
          5996 => x"44",
          5997 => x"76",
          5998 => x"81",
          5999 => x"38",
          6000 => x"ff",
          6001 => x"83",
          6002 => x"fd",
          6003 => x"1a",
          6004 => x"f8",
          6005 => x"e7",
          6006 => x"31",
          6007 => x"f8",
          6008 => x"90",
          6009 => x"58",
          6010 => x"26",
          6011 => x"80",
          6012 => x"05",
          6013 => x"f8",
          6014 => x"70",
          6015 => x"34",
          6016 => x"f4",
          6017 => x"76",
          6018 => x"58",
          6019 => x"90",
          6020 => x"81",
          6021 => x"79",
          6022 => x"38",
          6023 => x"79",
          6024 => x"75",
          6025 => x"23",
          6026 => x"80",
          6027 => x"94",
          6028 => x"39",
          6029 => x"92",
          6030 => x"39",
          6031 => x"f8",
          6032 => x"8e",
          6033 => x"83",
          6034 => x"f1",
          6035 => x"f8",
          6036 => x"5a",
          6037 => x"1a",
          6038 => x"80",
          6039 => x"e9",
          6040 => x"39",
          6041 => x"02",
          6042 => x"84",
          6043 => x"54",
          6044 => x"2e",
          6045 => x"51",
          6046 => x"80",
          6047 => x"e4",
          6048 => x"0d",
          6049 => x"73",
          6050 => x"3f",
          6051 => x"b8",
          6052 => x"3d",
          6053 => x"3d",
          6054 => x"05",
          6055 => x"0b",
          6056 => x"33",
          6057 => x"06",
          6058 => x"11",
          6059 => x"55",
          6060 => x"2e",
          6061 => x"81",
          6062 => x"83",
          6063 => x"74",
          6064 => x"b8",
          6065 => x"3d",
          6066 => x"f6",
          6067 => x"82",
          6068 => x"2e",
          6069 => x"73",
          6070 => x"71",
          6071 => x"70",
          6072 => x"5d",
          6073 => x"83",
          6074 => x"ff",
          6075 => x"7b",
          6076 => x"81",
          6077 => x"7b",
          6078 => x"32",
          6079 => x"80",
          6080 => x"5c",
          6081 => x"80",
          6082 => x"38",
          6083 => x"33",
          6084 => x"33",
          6085 => x"33",
          6086 => x"12",
          6087 => x"80",
          6088 => x"92",
          6089 => x"5d",
          6090 => x"05",
          6091 => x"ff",
          6092 => x"e9",
          6093 => x"55",
          6094 => x"2e",
          6095 => x"81",
          6096 => x"86",
          6097 => x"34",
          6098 => x"c0",
          6099 => x"87",
          6100 => x"08",
          6101 => x"2e",
          6102 => x"ee",
          6103 => x"57",
          6104 => x"94",
          6105 => x"14",
          6106 => x"06",
          6107 => x"f9",
          6108 => x"38",
          6109 => x"f6",
          6110 => x"70",
          6111 => x"83",
          6112 => x"33",
          6113 => x"72",
          6114 => x"c1",
          6115 => x"ff",
          6116 => x"38",
          6117 => x"98",
          6118 => x"81",
          6119 => x"79",
          6120 => x"85",
          6121 => x"83",
          6122 => x"34",
          6123 => x"14",
          6124 => x"8e",
          6125 => x"14",
          6126 => x"06",
          6127 => x"74",
          6128 => x"38",
          6129 => x"33",
          6130 => x"70",
          6131 => x"56",
          6132 => x"f6",
          6133 => x"81",
          6134 => x"86",
          6135 => x"70",
          6136 => x"54",
          6137 => x"2e",
          6138 => x"81",
          6139 => x"bd",
          6140 => x"81",
          6141 => x"80",
          6142 => x"38",
          6143 => x"f6",
          6144 => x"0b",
          6145 => x"33",
          6146 => x"08",
          6147 => x"33",
          6148 => x"c0",
          6149 => x"bf",
          6150 => x"42",
          6151 => x"56",
          6152 => x"16",
          6153 => x"81",
          6154 => x"38",
          6155 => x"16",
          6156 => x"80",
          6157 => x"38",
          6158 => x"16",
          6159 => x"81",
          6160 => x"38",
          6161 => x"16",
          6162 => x"81",
          6163 => x"81",
          6164 => x"73",
          6165 => x"8d",
          6166 => x"ac",
          6167 => x"72",
          6168 => x"da",
          6169 => x"ff",
          6170 => x"81",
          6171 => x"8c",
          6172 => x"ac",
          6173 => x"81",
          6174 => x"80",
          6175 => x"b8",
          6176 => x"05",
          6177 => x"9c",
          6178 => x"73",
          6179 => x"ec",
          6180 => x"87",
          6181 => x"08",
          6182 => x"0c",
          6183 => x"70",
          6184 => x"57",
          6185 => x"27",
          6186 => x"76",
          6187 => x"34",
          6188 => x"c0",
          6189 => x"19",
          6190 => x"26",
          6191 => x"72",
          6192 => x"c8",
          6193 => x"79",
          6194 => x"f6",
          6195 => x"73",
          6196 => x"38",
          6197 => x"87",
          6198 => x"08",
          6199 => x"7d",
          6200 => x"38",
          6201 => x"f6",
          6202 => x"54",
          6203 => x"83",
          6204 => x"73",
          6205 => x"34",
          6206 => x"9c",
          6207 => x"ec",
          6208 => x"ff",
          6209 => x"81",
          6210 => x"83",
          6211 => x"33",
          6212 => x"e0",
          6213 => x"34",
          6214 => x"fc",
          6215 => x"f6",
          6216 => x"72",
          6217 => x"9c",
          6218 => x"2e",
          6219 => x"80",
          6220 => x"81",
          6221 => x"8a",
          6222 => x"fe",
          6223 => x"74",
          6224 => x"59",
          6225 => x"9b",
          6226 => x"2e",
          6227 => x"83",
          6228 => x"81",
          6229 => x"38",
          6230 => x"80",
          6231 => x"81",
          6232 => x"87",
          6233 => x"98",
          6234 => x"72",
          6235 => x"38",
          6236 => x"9c",
          6237 => x"70",
          6238 => x"76",
          6239 => x"06",
          6240 => x"71",
          6241 => x"53",
          6242 => x"80",
          6243 => x"38",
          6244 => x"10",
          6245 => x"76",
          6246 => x"78",
          6247 => x"f4",
          6248 => x"5b",
          6249 => x"87",
          6250 => x"08",
          6251 => x"0c",
          6252 => x"39",
          6253 => x"81",
          6254 => x"38",
          6255 => x"06",
          6256 => x"39",
          6257 => x"9b",
          6258 => x"2e",
          6259 => x"80",
          6260 => x"da",
          6261 => x"72",
          6262 => x"e8",
          6263 => x"32",
          6264 => x"80",
          6265 => x"40",
          6266 => x"8a",
          6267 => x"2e",
          6268 => x"f9",
          6269 => x"ff",
          6270 => x"38",
          6271 => x"10",
          6272 => x"f6",
          6273 => x"33",
          6274 => x"7c",
          6275 => x"38",
          6276 => x"81",
          6277 => x"57",
          6278 => x"e2",
          6279 => x"db",
          6280 => x"80",
          6281 => x"38",
          6282 => x"33",
          6283 => x"91",
          6284 => x"ff",
          6285 => x"51",
          6286 => x"78",
          6287 => x"0c",
          6288 => x"04",
          6289 => x"81",
          6290 => x"f6",
          6291 => x"ff",
          6292 => x"83",
          6293 => x"33",
          6294 => x"7a",
          6295 => x"15",
          6296 => x"39",
          6297 => x"f6",
          6298 => x"ff",
          6299 => x"98",
          6300 => x"0b",
          6301 => x"15",
          6302 => x"39",
          6303 => x"06",
          6304 => x"ff",
          6305 => x"38",
          6306 => x"16",
          6307 => x"75",
          6308 => x"38",
          6309 => x"06",
          6310 => x"2e",
          6311 => x"fb",
          6312 => x"f6",
          6313 => x"fa",
          6314 => x"98",
          6315 => x"55",
          6316 => x"fb",
          6317 => x"c0",
          6318 => x"83",
          6319 => x"76",
          6320 => x"59",
          6321 => x"ff",
          6322 => x"98",
          6323 => x"ca",
          6324 => x"f6",
          6325 => x"09",
          6326 => x"72",
          6327 => x"72",
          6328 => x"34",
          6329 => x"f6",
          6330 => x"f6",
          6331 => x"f6",
          6332 => x"83",
          6333 => x"83",
          6334 => x"5d",
          6335 => x"5c",
          6336 => x"9c",
          6337 => x"2e",
          6338 => x"fc",
          6339 => x"59",
          6340 => x"fc",
          6341 => x"81",
          6342 => x"06",
          6343 => x"fd",
          6344 => x"76",
          6345 => x"54",
          6346 => x"80",
          6347 => x"db",
          6348 => x"75",
          6349 => x"54",
          6350 => x"db",
          6351 => x"f7",
          6352 => x"0b",
          6353 => x"33",
          6354 => x"83",
          6355 => x"73",
          6356 => x"34",
          6357 => x"95",
          6358 => x"83",
          6359 => x"84",
          6360 => x"38",
          6361 => x"f6",
          6362 => x"ff",
          6363 => x"d7",
          6364 => x"ff",
          6365 => x"57",
          6366 => x"79",
          6367 => x"80",
          6368 => x"f8",
          6369 => x"81",
          6370 => x"15",
          6371 => x"73",
          6372 => x"80",
          6373 => x"f8",
          6374 => x"b6",
          6375 => x"81",
          6376 => x"ff",
          6377 => x"75",
          6378 => x"80",
          6379 => x"f8",
          6380 => x"59",
          6381 => x"81",
          6382 => x"ff",
          6383 => x"ff",
          6384 => x"39",
          6385 => x"95",
          6386 => x"08",
          6387 => x"c8",
          6388 => x"f6",
          6389 => x"83",
          6390 => x"83",
          6391 => x"59",
          6392 => x"80",
          6393 => x"51",
          6394 => x"82",
          6395 => x"fa",
          6396 => x"0b",
          6397 => x"08",
          6398 => x"a3",
          6399 => x"13",
          6400 => x"f0",
          6401 => x"e0",
          6402 => x"0b",
          6403 => x"08",
          6404 => x"0b",
          6405 => x"80",
          6406 => x"80",
          6407 => x"c0",
          6408 => x"83",
          6409 => x"55",
          6410 => x"05",
          6411 => x"98",
          6412 => x"87",
          6413 => x"08",
          6414 => x"2e",
          6415 => x"14",
          6416 => x"98",
          6417 => x"52",
          6418 => x"87",
          6419 => x"fe",
          6420 => x"87",
          6421 => x"08",
          6422 => x"70",
          6423 => x"c8",
          6424 => x"71",
          6425 => x"c0",
          6426 => x"98",
          6427 => x"ce",
          6428 => x"87",
          6429 => x"08",
          6430 => x"98",
          6431 => x"74",
          6432 => x"38",
          6433 => x"87",
          6434 => x"08",
          6435 => x"73",
          6436 => x"71",
          6437 => x"db",
          6438 => x"98",
          6439 => x"72",
          6440 => x"38",
          6441 => x"55",
          6442 => x"81",
          6443 => x"53",
          6444 => x"98",
          6445 => x"ff",
          6446 => x"fe",
          6447 => x"ff",
          6448 => x"76",
          6449 => x"0c",
          6450 => x"04",
          6451 => x"b8",
          6452 => x"3d",
          6453 => x"3d",
          6454 => x"84",
          6455 => x"33",
          6456 => x"0b",
          6457 => x"08",
          6458 => x"87",
          6459 => x"06",
          6460 => x"2a",
          6461 => x"55",
          6462 => x"15",
          6463 => x"2a",
          6464 => x"15",
          6465 => x"2a",
          6466 => x"15",
          6467 => x"15",
          6468 => x"f0",
          6469 => x"82",
          6470 => x"f2",
          6471 => x"80",
          6472 => x"85",
          6473 => x"f0",
          6474 => x"fe",
          6475 => x"34",
          6476 => x"f0",
          6477 => x"87",
          6478 => x"08",
          6479 => x"08",
          6480 => x"90",
          6481 => x"c0",
          6482 => x"52",
          6483 => x"9c",
          6484 => x"72",
          6485 => x"81",
          6486 => x"c0",
          6487 => x"56",
          6488 => x"27",
          6489 => x"81",
          6490 => x"38",
          6491 => x"a4",
          6492 => x"55",
          6493 => x"80",
          6494 => x"55",
          6495 => x"80",
          6496 => x"c0",
          6497 => x"80",
          6498 => x"53",
          6499 => x"9c",
          6500 => x"c0",
          6501 => x"55",
          6502 => x"f6",
          6503 => x"33",
          6504 => x"9c",
          6505 => x"70",
          6506 => x"38",
          6507 => x"2e",
          6508 => x"c0",
          6509 => x"55",
          6510 => x"83",
          6511 => x"71",
          6512 => x"70",
          6513 => x"57",
          6514 => x"2e",
          6515 => x"74",
          6516 => x"52",
          6517 => x"38",
          6518 => x"81",
          6519 => x"75",
          6520 => x"c6",
          6521 => x"80",
          6522 => x"52",
          6523 => x"92",
          6524 => x"81",
          6525 => x"71",
          6526 => x"53",
          6527 => x"26",
          6528 => x"84",
          6529 => x"88",
          6530 => x"81",
          6531 => x"e4",
          6532 => x"0d",
          6533 => x"c2",
          6534 => x"0d",
          6535 => x"05",
          6536 => x"56",
          6537 => x"83",
          6538 => x"77",
          6539 => x"fc",
          6540 => x"70",
          6541 => x"07",
          6542 => x"57",
          6543 => x"34",
          6544 => x"51",
          6545 => x"34",
          6546 => x"52",
          6547 => x"34",
          6548 => x"34",
          6549 => x"f0",
          6550 => x"11",
          6551 => x"56",
          6552 => x"70",
          6553 => x"38",
          6554 => x"05",
          6555 => x"70",
          6556 => x"34",
          6557 => x"f0",
          6558 => x"f0",
          6559 => x"82",
          6560 => x"f2",
          6561 => x"80",
          6562 => x"85",
          6563 => x"f0",
          6564 => x"fe",
          6565 => x"34",
          6566 => x"f0",
          6567 => x"87",
          6568 => x"08",
          6569 => x"08",
          6570 => x"90",
          6571 => x"c0",
          6572 => x"52",
          6573 => x"9c",
          6574 => x"72",
          6575 => x"81",
          6576 => x"c0",
          6577 => x"56",
          6578 => x"27",
          6579 => x"81",
          6580 => x"38",
          6581 => x"a4",
          6582 => x"55",
          6583 => x"80",
          6584 => x"55",
          6585 => x"80",
          6586 => x"c0",
          6587 => x"80",
          6588 => x"53",
          6589 => x"9c",
          6590 => x"c0",
          6591 => x"55",
          6592 => x"f6",
          6593 => x"33",
          6594 => x"9c",
          6595 => x"70",
          6596 => x"38",
          6597 => x"2e",
          6598 => x"c0",
          6599 => x"55",
          6600 => x"83",
          6601 => x"71",
          6602 => x"70",
          6603 => x"57",
          6604 => x"2e",
          6605 => x"81",
          6606 => x"71",
          6607 => x"74",
          6608 => x"ff",
          6609 => x"80",
          6610 => x"81",
          6611 => x"b8",
          6612 => x"3d",
          6613 => x"51",
          6614 => x"3d",
          6615 => x"f0",
          6616 => x"d0",
          6617 => x"0b",
          6618 => x"08",
          6619 => x"0b",
          6620 => x"80",
          6621 => x"80",
          6622 => x"c0",
          6623 => x"83",
          6624 => x"56",
          6625 => x"05",
          6626 => x"98",
          6627 => x"87",
          6628 => x"08",
          6629 => x"2e",
          6630 => x"15",
          6631 => x"98",
          6632 => x"52",
          6633 => x"87",
          6634 => x"fe",
          6635 => x"87",
          6636 => x"08",
          6637 => x"70",
          6638 => x"c8",
          6639 => x"71",
          6640 => x"c0",
          6641 => x"98",
          6642 => x"ce",
          6643 => x"87",
          6644 => x"08",
          6645 => x"98",
          6646 => x"70",
          6647 => x"38",
          6648 => x"87",
          6649 => x"08",
          6650 => x"73",
          6651 => x"71",
          6652 => x"db",
          6653 => x"98",
          6654 => x"72",
          6655 => x"38",
          6656 => x"53",
          6657 => x"81",
          6658 => x"52",
          6659 => x"8a",
          6660 => x"ff",
          6661 => x"fe",
          6662 => x"39",
          6663 => x"83",
          6664 => x"fe",
          6665 => x"82",
          6666 => x"f9",
          6667 => x"b8",
          6668 => x"71",
          6669 => x"70",
          6670 => x"06",
          6671 => x"73",
          6672 => x"81",
          6673 => x"8b",
          6674 => x"2b",
          6675 => x"70",
          6676 => x"33",
          6677 => x"71",
          6678 => x"5c",
          6679 => x"53",
          6680 => x"52",
          6681 => x"80",
          6682 => x"af",
          6683 => x"82",
          6684 => x"12",
          6685 => x"2b",
          6686 => x"07",
          6687 => x"33",
          6688 => x"71",
          6689 => x"90",
          6690 => x"53",
          6691 => x"56",
          6692 => x"24",
          6693 => x"84",
          6694 => x"14",
          6695 => x"2b",
          6696 => x"07",
          6697 => x"88",
          6698 => x"56",
          6699 => x"13",
          6700 => x"ff",
          6701 => x"87",
          6702 => x"b8",
          6703 => x"17",
          6704 => x"85",
          6705 => x"88",
          6706 => x"88",
          6707 => x"59",
          6708 => x"84",
          6709 => x"85",
          6710 => x"b8",
          6711 => x"52",
          6712 => x"13",
          6713 => x"87",
          6714 => x"b8",
          6715 => x"74",
          6716 => x"73",
          6717 => x"84",
          6718 => x"16",
          6719 => x"12",
          6720 => x"2b",
          6721 => x"80",
          6722 => x"2a",
          6723 => x"52",
          6724 => x"75",
          6725 => x"89",
          6726 => x"86",
          6727 => x"13",
          6728 => x"2b",
          6729 => x"07",
          6730 => x"16",
          6731 => x"33",
          6732 => x"07",
          6733 => x"58",
          6734 => x"53",
          6735 => x"84",
          6736 => x"85",
          6737 => x"b8",
          6738 => x"16",
          6739 => x"85",
          6740 => x"8b",
          6741 => x"2b",
          6742 => x"5a",
          6743 => x"86",
          6744 => x"13",
          6745 => x"2b",
          6746 => x"2a",
          6747 => x"52",
          6748 => x"34",
          6749 => x"34",
          6750 => x"08",
          6751 => x"81",
          6752 => x"88",
          6753 => x"ff",
          6754 => x"88",
          6755 => x"54",
          6756 => x"34",
          6757 => x"34",
          6758 => x"08",
          6759 => x"33",
          6760 => x"71",
          6761 => x"83",
          6762 => x"05",
          6763 => x"12",
          6764 => x"2b",
          6765 => x"2b",
          6766 => x"06",
          6767 => x"88",
          6768 => x"53",
          6769 => x"57",
          6770 => x"82",
          6771 => x"83",
          6772 => x"b8",
          6773 => x"17",
          6774 => x"12",
          6775 => x"2b",
          6776 => x"07",
          6777 => x"33",
          6778 => x"71",
          6779 => x"81",
          6780 => x"70",
          6781 => x"52",
          6782 => x"57",
          6783 => x"73",
          6784 => x"14",
          6785 => x"d4",
          6786 => x"82",
          6787 => x"12",
          6788 => x"2b",
          6789 => x"07",
          6790 => x"33",
          6791 => x"71",
          6792 => x"90",
          6793 => x"53",
          6794 => x"57",
          6795 => x"80",
          6796 => x"38",
          6797 => x"13",
          6798 => x"2b",
          6799 => x"80",
          6800 => x"2a",
          6801 => x"76",
          6802 => x"81",
          6803 => x"b8",
          6804 => x"17",
          6805 => x"12",
          6806 => x"2b",
          6807 => x"07",
          6808 => x"14",
          6809 => x"33",
          6810 => x"07",
          6811 => x"57",
          6812 => x"58",
          6813 => x"72",
          6814 => x"75",
          6815 => x"89",
          6816 => x"f9",
          6817 => x"84",
          6818 => x"58",
          6819 => x"2e",
          6820 => x"80",
          6821 => x"77",
          6822 => x"3f",
          6823 => x"04",
          6824 => x"0b",
          6825 => x"0c",
          6826 => x"84",
          6827 => x"82",
          6828 => x"76",
          6829 => x"f4",
          6830 => x"c6",
          6831 => x"d4",
          6832 => x"75",
          6833 => x"81",
          6834 => x"b8",
          6835 => x"76",
          6836 => x"81",
          6837 => x"34",
          6838 => x"08",
          6839 => x"17",
          6840 => x"87",
          6841 => x"b8",
          6842 => x"b8",
          6843 => x"05",
          6844 => x"07",
          6845 => x"ff",
          6846 => x"2a",
          6847 => x"56",
          6848 => x"34",
          6849 => x"34",
          6850 => x"22",
          6851 => x"10",
          6852 => x"08",
          6853 => x"55",
          6854 => x"15",
          6855 => x"83",
          6856 => x"ee",
          6857 => x"0d",
          6858 => x"53",
          6859 => x"72",
          6860 => x"fb",
          6861 => x"82",
          6862 => x"ff",
          6863 => x"51",
          6864 => x"ff",
          6865 => x"d4",
          6866 => x"33",
          6867 => x"71",
          6868 => x"70",
          6869 => x"58",
          6870 => x"ff",
          6871 => x"2e",
          6872 => x"75",
          6873 => x"17",
          6874 => x"12",
          6875 => x"2b",
          6876 => x"ff",
          6877 => x"31",
          6878 => x"ff",
          6879 => x"27",
          6880 => x"5c",
          6881 => x"74",
          6882 => x"70",
          6883 => x"38",
          6884 => x"58",
          6885 => x"85",
          6886 => x"88",
          6887 => x"5a",
          6888 => x"73",
          6889 => x"2e",
          6890 => x"74",
          6891 => x"76",
          6892 => x"11",
          6893 => x"12",
          6894 => x"2b",
          6895 => x"ff",
          6896 => x"56",
          6897 => x"59",
          6898 => x"83",
          6899 => x"80",
          6900 => x"26",
          6901 => x"78",
          6902 => x"2e",
          6903 => x"72",
          6904 => x"88",
          6905 => x"70",
          6906 => x"11",
          6907 => x"80",
          6908 => x"2a",
          6909 => x"56",
          6910 => x"34",
          6911 => x"34",
          6912 => x"08",
          6913 => x"2a",
          6914 => x"82",
          6915 => x"83",
          6916 => x"b8",
          6917 => x"19",
          6918 => x"12",
          6919 => x"2b",
          6920 => x"2b",
          6921 => x"06",
          6922 => x"83",
          6923 => x"70",
          6924 => x"58",
          6925 => x"52",
          6926 => x"12",
          6927 => x"ff",
          6928 => x"83",
          6929 => x"b8",
          6930 => x"54",
          6931 => x"72",
          6932 => x"84",
          6933 => x"70",
          6934 => x"33",
          6935 => x"71",
          6936 => x"83",
          6937 => x"05",
          6938 => x"53",
          6939 => x"15",
          6940 => x"15",
          6941 => x"d4",
          6942 => x"55",
          6943 => x"11",
          6944 => x"33",
          6945 => x"07",
          6946 => x"54",
          6947 => x"70",
          6948 => x"71",
          6949 => x"84",
          6950 => x"70",
          6951 => x"33",
          6952 => x"71",
          6953 => x"83",
          6954 => x"05",
          6955 => x"5a",
          6956 => x"15",
          6957 => x"15",
          6958 => x"d4",
          6959 => x"55",
          6960 => x"11",
          6961 => x"33",
          6962 => x"07",
          6963 => x"54",
          6964 => x"70",
          6965 => x"79",
          6966 => x"84",
          6967 => x"18",
          6968 => x"70",
          6969 => x"0c",
          6970 => x"04",
          6971 => x"87",
          6972 => x"8b",
          6973 => x"2b",
          6974 => x"84",
          6975 => x"18",
          6976 => x"2b",
          6977 => x"2a",
          6978 => x"53",
          6979 => x"84",
          6980 => x"85",
          6981 => x"b8",
          6982 => x"19",
          6983 => x"85",
          6984 => x"8b",
          6985 => x"2b",
          6986 => x"86",
          6987 => x"15",
          6988 => x"2b",
          6989 => x"2a",
          6990 => x"52",
          6991 => x"52",
          6992 => x"34",
          6993 => x"34",
          6994 => x"08",
          6995 => x"81",
          6996 => x"88",
          6997 => x"ff",
          6998 => x"88",
          6999 => x"54",
          7000 => x"34",
          7001 => x"34",
          7002 => x"08",
          7003 => x"51",
          7004 => x"f9",
          7005 => x"84",
          7006 => x"58",
          7007 => x"2e",
          7008 => x"54",
          7009 => x"73",
          7010 => x"0c",
          7011 => x"04",
          7012 => x"91",
          7013 => x"e4",
          7014 => x"e4",
          7015 => x"0d",
          7016 => x"f4",
          7017 => x"d4",
          7018 => x"0b",
          7019 => x"23",
          7020 => x"53",
          7021 => x"ff",
          7022 => x"cd",
          7023 => x"b8",
          7024 => x"76",
          7025 => x"0b",
          7026 => x"84",
          7027 => x"54",
          7028 => x"34",
          7029 => x"15",
          7030 => x"d4",
          7031 => x"86",
          7032 => x"0b",
          7033 => x"84",
          7034 => x"84",
          7035 => x"ff",
          7036 => x"80",
          7037 => x"ff",
          7038 => x"88",
          7039 => x"55",
          7040 => x"17",
          7041 => x"17",
          7042 => x"d0",
          7043 => x"10",
          7044 => x"d4",
          7045 => x"05",
          7046 => x"82",
          7047 => x"0b",
          7048 => x"77",
          7049 => x"2e",
          7050 => x"fe",
          7051 => x"3d",
          7052 => x"41",
          7053 => x"84",
          7054 => x"59",
          7055 => x"61",
          7056 => x"38",
          7057 => x"85",
          7058 => x"80",
          7059 => x"38",
          7060 => x"60",
          7061 => x"7f",
          7062 => x"2a",
          7063 => x"83",
          7064 => x"55",
          7065 => x"ff",
          7066 => x"78",
          7067 => x"70",
          7068 => x"06",
          7069 => x"7a",
          7070 => x"81",
          7071 => x"88",
          7072 => x"75",
          7073 => x"ff",
          7074 => x"10",
          7075 => x"05",
          7076 => x"61",
          7077 => x"81",
          7078 => x"88",
          7079 => x"90",
          7080 => x"2c",
          7081 => x"46",
          7082 => x"43",
          7083 => x"59",
          7084 => x"42",
          7085 => x"85",
          7086 => x"15",
          7087 => x"33",
          7088 => x"07",
          7089 => x"10",
          7090 => x"81",
          7091 => x"98",
          7092 => x"2b",
          7093 => x"53",
          7094 => x"80",
          7095 => x"c9",
          7096 => x"27",
          7097 => x"63",
          7098 => x"62",
          7099 => x"38",
          7100 => x"85",
          7101 => x"1b",
          7102 => x"25",
          7103 => x"63",
          7104 => x"79",
          7105 => x"38",
          7106 => x"33",
          7107 => x"71",
          7108 => x"83",
          7109 => x"11",
          7110 => x"12",
          7111 => x"2b",
          7112 => x"07",
          7113 => x"52",
          7114 => x"58",
          7115 => x"8c",
          7116 => x"1e",
          7117 => x"83",
          7118 => x"8b",
          7119 => x"2b",
          7120 => x"86",
          7121 => x"12",
          7122 => x"2b",
          7123 => x"07",
          7124 => x"14",
          7125 => x"33",
          7126 => x"07",
          7127 => x"59",
          7128 => x"5b",
          7129 => x"5c",
          7130 => x"84",
          7131 => x"85",
          7132 => x"b8",
          7133 => x"17",
          7134 => x"85",
          7135 => x"8b",
          7136 => x"2b",
          7137 => x"86",
          7138 => x"15",
          7139 => x"2b",
          7140 => x"2a",
          7141 => x"52",
          7142 => x"57",
          7143 => x"34",
          7144 => x"34",
          7145 => x"08",
          7146 => x"81",
          7147 => x"88",
          7148 => x"ff",
          7149 => x"88",
          7150 => x"5e",
          7151 => x"34",
          7152 => x"34",
          7153 => x"08",
          7154 => x"11",
          7155 => x"33",
          7156 => x"71",
          7157 => x"74",
          7158 => x"81",
          7159 => x"88",
          7160 => x"88",
          7161 => x"45",
          7162 => x"55",
          7163 => x"34",
          7164 => x"34",
          7165 => x"08",
          7166 => x"33",
          7167 => x"71",
          7168 => x"83",
          7169 => x"05",
          7170 => x"83",
          7171 => x"88",
          7172 => x"88",
          7173 => x"45",
          7174 => x"55",
          7175 => x"1a",
          7176 => x"1a",
          7177 => x"d4",
          7178 => x"82",
          7179 => x"12",
          7180 => x"2b",
          7181 => x"62",
          7182 => x"2b",
          7183 => x"5d",
          7184 => x"05",
          7185 => x"fd",
          7186 => x"d4",
          7187 => x"05",
          7188 => x"1c",
          7189 => x"ff",
          7190 => x"5f",
          7191 => x"81",
          7192 => x"54",
          7193 => x"e4",
          7194 => x"0d",
          7195 => x"f4",
          7196 => x"d4",
          7197 => x"0b",
          7198 => x"23",
          7199 => x"53",
          7200 => x"ff",
          7201 => x"c7",
          7202 => x"b8",
          7203 => x"60",
          7204 => x"0b",
          7205 => x"84",
          7206 => x"5d",
          7207 => x"34",
          7208 => x"1e",
          7209 => x"d4",
          7210 => x"86",
          7211 => x"0b",
          7212 => x"84",
          7213 => x"84",
          7214 => x"ff",
          7215 => x"80",
          7216 => x"ff",
          7217 => x"88",
          7218 => x"5b",
          7219 => x"18",
          7220 => x"18",
          7221 => x"d0",
          7222 => x"10",
          7223 => x"d4",
          7224 => x"05",
          7225 => x"82",
          7226 => x"0b",
          7227 => x"84",
          7228 => x"57",
          7229 => x"38",
          7230 => x"82",
          7231 => x"54",
          7232 => x"fe",
          7233 => x"51",
          7234 => x"84",
          7235 => x"84",
          7236 => x"95",
          7237 => x"61",
          7238 => x"d4",
          7239 => x"2b",
          7240 => x"44",
          7241 => x"33",
          7242 => x"71",
          7243 => x"81",
          7244 => x"70",
          7245 => x"44",
          7246 => x"63",
          7247 => x"81",
          7248 => x"84",
          7249 => x"05",
          7250 => x"57",
          7251 => x"19",
          7252 => x"19",
          7253 => x"d4",
          7254 => x"70",
          7255 => x"33",
          7256 => x"07",
          7257 => x"8f",
          7258 => x"74",
          7259 => x"ff",
          7260 => x"88",
          7261 => x"47",
          7262 => x"5d",
          7263 => x"05",
          7264 => x"ff",
          7265 => x"63",
          7266 => x"84",
          7267 => x"1e",
          7268 => x"34",
          7269 => x"34",
          7270 => x"d4",
          7271 => x"05",
          7272 => x"3f",
          7273 => x"bc",
          7274 => x"31",
          7275 => x"ff",
          7276 => x"fa",
          7277 => x"81",
          7278 => x"76",
          7279 => x"ff",
          7280 => x"17",
          7281 => x"33",
          7282 => x"07",
          7283 => x"10",
          7284 => x"81",
          7285 => x"98",
          7286 => x"2b",
          7287 => x"53",
          7288 => x"45",
          7289 => x"25",
          7290 => x"ff",
          7291 => x"78",
          7292 => x"38",
          7293 => x"8b",
          7294 => x"83",
          7295 => x"5b",
          7296 => x"fc",
          7297 => x"8f",
          7298 => x"f4",
          7299 => x"d4",
          7300 => x"0b",
          7301 => x"23",
          7302 => x"53",
          7303 => x"ff",
          7304 => x"c4",
          7305 => x"b8",
          7306 => x"7e",
          7307 => x"0b",
          7308 => x"84",
          7309 => x"59",
          7310 => x"34",
          7311 => x"1a",
          7312 => x"d4",
          7313 => x"86",
          7314 => x"0b",
          7315 => x"84",
          7316 => x"84",
          7317 => x"ff",
          7318 => x"80",
          7319 => x"ff",
          7320 => x"88",
          7321 => x"57",
          7322 => x"88",
          7323 => x"64",
          7324 => x"84",
          7325 => x"70",
          7326 => x"84",
          7327 => x"05",
          7328 => x"43",
          7329 => x"05",
          7330 => x"83",
          7331 => x"ee",
          7332 => x"24",
          7333 => x"61",
          7334 => x"06",
          7335 => x"27",
          7336 => x"fc",
          7337 => x"80",
          7338 => x"38",
          7339 => x"fb",
          7340 => x"73",
          7341 => x"0c",
          7342 => x"04",
          7343 => x"11",
          7344 => x"33",
          7345 => x"71",
          7346 => x"7a",
          7347 => x"33",
          7348 => x"71",
          7349 => x"83",
          7350 => x"05",
          7351 => x"85",
          7352 => x"88",
          7353 => x"88",
          7354 => x"45",
          7355 => x"58",
          7356 => x"56",
          7357 => x"05",
          7358 => x"85",
          7359 => x"b8",
          7360 => x"17",
          7361 => x"85",
          7362 => x"8b",
          7363 => x"2b",
          7364 => x"86",
          7365 => x"15",
          7366 => x"2b",
          7367 => x"2a",
          7368 => x"48",
          7369 => x"41",
          7370 => x"05",
          7371 => x"87",
          7372 => x"b8",
          7373 => x"70",
          7374 => x"33",
          7375 => x"07",
          7376 => x"06",
          7377 => x"5f",
          7378 => x"7b",
          7379 => x"81",
          7380 => x"b8",
          7381 => x"1f",
          7382 => x"83",
          7383 => x"8b",
          7384 => x"2b",
          7385 => x"73",
          7386 => x"33",
          7387 => x"07",
          7388 => x"5e",
          7389 => x"43",
          7390 => x"76",
          7391 => x"81",
          7392 => x"b8",
          7393 => x"1f",
          7394 => x"12",
          7395 => x"2b",
          7396 => x"07",
          7397 => x"14",
          7398 => x"33",
          7399 => x"07",
          7400 => x"40",
          7401 => x"40",
          7402 => x"78",
          7403 => x"60",
          7404 => x"84",
          7405 => x"70",
          7406 => x"33",
          7407 => x"71",
          7408 => x"66",
          7409 => x"70",
          7410 => x"52",
          7411 => x"05",
          7412 => x"fe",
          7413 => x"84",
          7414 => x"1e",
          7415 => x"83",
          7416 => x"5c",
          7417 => x"39",
          7418 => x"0b",
          7419 => x"0c",
          7420 => x"84",
          7421 => x"82",
          7422 => x"7f",
          7423 => x"f4",
          7424 => x"fe",
          7425 => x"d4",
          7426 => x"76",
          7427 => x"81",
          7428 => x"b8",
          7429 => x"7f",
          7430 => x"81",
          7431 => x"34",
          7432 => x"08",
          7433 => x"15",
          7434 => x"87",
          7435 => x"b8",
          7436 => x"b8",
          7437 => x"05",
          7438 => x"07",
          7439 => x"ff",
          7440 => x"2a",
          7441 => x"5e",
          7442 => x"34",
          7443 => x"34",
          7444 => x"22",
          7445 => x"10",
          7446 => x"08",
          7447 => x"5c",
          7448 => x"1c",
          7449 => x"83",
          7450 => x"51",
          7451 => x"7f",
          7452 => x"39",
          7453 => x"87",
          7454 => x"8b",
          7455 => x"2b",
          7456 => x"84",
          7457 => x"1d",
          7458 => x"2b",
          7459 => x"2a",
          7460 => x"43",
          7461 => x"61",
          7462 => x"63",
          7463 => x"34",
          7464 => x"08",
          7465 => x"11",
          7466 => x"33",
          7467 => x"71",
          7468 => x"74",
          7469 => x"33",
          7470 => x"71",
          7471 => x"70",
          7472 => x"5f",
          7473 => x"56",
          7474 => x"64",
          7475 => x"78",
          7476 => x"34",
          7477 => x"08",
          7478 => x"81",
          7479 => x"88",
          7480 => x"ff",
          7481 => x"88",
          7482 => x"58",
          7483 => x"34",
          7484 => x"34",
          7485 => x"08",
          7486 => x"33",
          7487 => x"71",
          7488 => x"83",
          7489 => x"05",
          7490 => x"12",
          7491 => x"2b",
          7492 => x"2b",
          7493 => x"06",
          7494 => x"88",
          7495 => x"5d",
          7496 => x"5d",
          7497 => x"82",
          7498 => x"83",
          7499 => x"b8",
          7500 => x"1f",
          7501 => x"12",
          7502 => x"2b",
          7503 => x"07",
          7504 => x"33",
          7505 => x"71",
          7506 => x"81",
          7507 => x"70",
          7508 => x"5d",
          7509 => x"5a",
          7510 => x"60",
          7511 => x"81",
          7512 => x"83",
          7513 => x"5b",
          7514 => x"86",
          7515 => x"16",
          7516 => x"2b",
          7517 => x"07",
          7518 => x"18",
          7519 => x"33",
          7520 => x"07",
          7521 => x"5e",
          7522 => x"41",
          7523 => x"1e",
          7524 => x"1e",
          7525 => x"d4",
          7526 => x"84",
          7527 => x"12",
          7528 => x"2b",
          7529 => x"07",
          7530 => x"14",
          7531 => x"33",
          7532 => x"07",
          7533 => x"44",
          7534 => x"5a",
          7535 => x"7c",
          7536 => x"34",
          7537 => x"05",
          7538 => x"d4",
          7539 => x"33",
          7540 => x"71",
          7541 => x"81",
          7542 => x"70",
          7543 => x"5b",
          7544 => x"75",
          7545 => x"16",
          7546 => x"d4",
          7547 => x"70",
          7548 => x"33",
          7549 => x"71",
          7550 => x"74",
          7551 => x"81",
          7552 => x"88",
          7553 => x"83",
          7554 => x"f8",
          7555 => x"63",
          7556 => x"54",
          7557 => x"59",
          7558 => x"7f",
          7559 => x"7b",
          7560 => x"84",
          7561 => x"70",
          7562 => x"81",
          7563 => x"8b",
          7564 => x"2b",
          7565 => x"70",
          7566 => x"33",
          7567 => x"07",
          7568 => x"06",
          7569 => x"5d",
          7570 => x"5b",
          7571 => x"75",
          7572 => x"81",
          7573 => x"b8",
          7574 => x"1f",
          7575 => x"83",
          7576 => x"8b",
          7577 => x"2b",
          7578 => x"86",
          7579 => x"12",
          7580 => x"2b",
          7581 => x"07",
          7582 => x"14",
          7583 => x"33",
          7584 => x"07",
          7585 => x"59",
          7586 => x"5c",
          7587 => x"5d",
          7588 => x"77",
          7589 => x"79",
          7590 => x"84",
          7591 => x"70",
          7592 => x"33",
          7593 => x"71",
          7594 => x"83",
          7595 => x"05",
          7596 => x"87",
          7597 => x"88",
          7598 => x"88",
          7599 => x"5e",
          7600 => x"41",
          7601 => x"16",
          7602 => x"16",
          7603 => x"d4",
          7604 => x"33",
          7605 => x"71",
          7606 => x"81",
          7607 => x"70",
          7608 => x"5c",
          7609 => x"79",
          7610 => x"1a",
          7611 => x"d4",
          7612 => x"82",
          7613 => x"12",
          7614 => x"2b",
          7615 => x"07",
          7616 => x"33",
          7617 => x"71",
          7618 => x"70",
          7619 => x"5c",
          7620 => x"5a",
          7621 => x"79",
          7622 => x"1a",
          7623 => x"d4",
          7624 => x"70",
          7625 => x"33",
          7626 => x"71",
          7627 => x"74",
          7628 => x"33",
          7629 => x"71",
          7630 => x"70",
          7631 => x"5c",
          7632 => x"5a",
          7633 => x"82",
          7634 => x"83",
          7635 => x"b8",
          7636 => x"1f",
          7637 => x"83",
          7638 => x"88",
          7639 => x"57",
          7640 => x"83",
          7641 => x"5a",
          7642 => x"84",
          7643 => x"b6",
          7644 => x"b8",
          7645 => x"84",
          7646 => x"05",
          7647 => x"ff",
          7648 => x"44",
          7649 => x"39",
          7650 => x"87",
          7651 => x"8b",
          7652 => x"2b",
          7653 => x"84",
          7654 => x"1d",
          7655 => x"2b",
          7656 => x"2a",
          7657 => x"43",
          7658 => x"61",
          7659 => x"63",
          7660 => x"34",
          7661 => x"08",
          7662 => x"11",
          7663 => x"33",
          7664 => x"71",
          7665 => x"74",
          7666 => x"33",
          7667 => x"71",
          7668 => x"70",
          7669 => x"41",
          7670 => x"59",
          7671 => x"64",
          7672 => x"7a",
          7673 => x"34",
          7674 => x"08",
          7675 => x"81",
          7676 => x"88",
          7677 => x"ff",
          7678 => x"88",
          7679 => x"42",
          7680 => x"34",
          7681 => x"34",
          7682 => x"08",
          7683 => x"33",
          7684 => x"71",
          7685 => x"83",
          7686 => x"05",
          7687 => x"12",
          7688 => x"2b",
          7689 => x"2b",
          7690 => x"06",
          7691 => x"88",
          7692 => x"5c",
          7693 => x"45",
          7694 => x"82",
          7695 => x"83",
          7696 => x"b8",
          7697 => x"1f",
          7698 => x"12",
          7699 => x"2b",
          7700 => x"07",
          7701 => x"33",
          7702 => x"71",
          7703 => x"81",
          7704 => x"70",
          7705 => x"5f",
          7706 => x"59",
          7707 => x"7d",
          7708 => x"1e",
          7709 => x"ff",
          7710 => x"f3",
          7711 => x"60",
          7712 => x"a1",
          7713 => x"e4",
          7714 => x"b8",
          7715 => x"2e",
          7716 => x"53",
          7717 => x"b8",
          7718 => x"fe",
          7719 => x"73",
          7720 => x"3f",
          7721 => x"7b",
          7722 => x"38",
          7723 => x"f9",
          7724 => x"7a",
          7725 => x"d4",
          7726 => x"76",
          7727 => x"38",
          7728 => x"8a",
          7729 => x"b8",
          7730 => x"3d",
          7731 => x"51",
          7732 => x"84",
          7733 => x"54",
          7734 => x"08",
          7735 => x"38",
          7736 => x"52",
          7737 => x"08",
          7738 => x"96",
          7739 => x"b8",
          7740 => x"3d",
          7741 => x"ff",
          7742 => x"b8",
          7743 => x"80",
          7744 => x"d0",
          7745 => x"80",
          7746 => x"84",
          7747 => x"fe",
          7748 => x"84",
          7749 => x"55",
          7750 => x"81",
          7751 => x"34",
          7752 => x"08",
          7753 => x"15",
          7754 => x"85",
          7755 => x"b8",
          7756 => x"76",
          7757 => x"81",
          7758 => x"34",
          7759 => x"08",
          7760 => x"22",
          7761 => x"80",
          7762 => x"83",
          7763 => x"70",
          7764 => x"51",
          7765 => x"88",
          7766 => x"89",
          7767 => x"b8",
          7768 => x"10",
          7769 => x"b8",
          7770 => x"f8",
          7771 => x"76",
          7772 => x"81",
          7773 => x"34",
          7774 => x"80",
          7775 => x"38",
          7776 => x"ff",
          7777 => x"8f",
          7778 => x"81",
          7779 => x"26",
          7780 => x"b8",
          7781 => x"52",
          7782 => x"e4",
          7783 => x"0d",
          7784 => x"0d",
          7785 => x"33",
          7786 => x"71",
          7787 => x"38",
          7788 => x"bb",
          7789 => x"e4",
          7790 => x"06",
          7791 => x"38",
          7792 => x"e0",
          7793 => x"b8",
          7794 => x"53",
          7795 => x"e4",
          7796 => x"0d",
          7797 => x"0d",
          7798 => x"02",
          7799 => x"05",
          7800 => x"57",
          7801 => x"76",
          7802 => x"38",
          7803 => x"17",
          7804 => x"81",
          7805 => x"55",
          7806 => x"73",
          7807 => x"87",
          7808 => x"0c",
          7809 => x"52",
          7810 => x"ca",
          7811 => x"e4",
          7812 => x"06",
          7813 => x"2e",
          7814 => x"c0",
          7815 => x"54",
          7816 => x"79",
          7817 => x"38",
          7818 => x"80",
          7819 => x"80",
          7820 => x"81",
          7821 => x"74",
          7822 => x"0c",
          7823 => x"04",
          7824 => x"81",
          7825 => x"ff",
          7826 => x"56",
          7827 => x"ff",
          7828 => x"39",
          7829 => x"7c",
          7830 => x"8c",
          7831 => x"33",
          7832 => x"59",
          7833 => x"74",
          7834 => x"84",
          7835 => x"33",
          7836 => x"06",
          7837 => x"73",
          7838 => x"58",
          7839 => x"c0",
          7840 => x"78",
          7841 => x"76",
          7842 => x"3f",
          7843 => x"08",
          7844 => x"55",
          7845 => x"a7",
          7846 => x"98",
          7847 => x"73",
          7848 => x"78",
          7849 => x"74",
          7850 => x"06",
          7851 => x"2e",
          7852 => x"54",
          7853 => x"84",
          7854 => x"8b",
          7855 => x"84",
          7856 => x"19",
          7857 => x"06",
          7858 => x"79",
          7859 => x"ac",
          7860 => x"fc",
          7861 => x"02",
          7862 => x"05",
          7863 => x"05",
          7864 => x"53",
          7865 => x"53",
          7866 => x"87",
          7867 => x"e0",
          7868 => x"72",
          7869 => x"83",
          7870 => x"38",
          7871 => x"c0",
          7872 => x"81",
          7873 => x"2e",
          7874 => x"71",
          7875 => x"70",
          7876 => x"38",
          7877 => x"84",
          7878 => x"86",
          7879 => x"88",
          7880 => x"0c",
          7881 => x"e4",
          7882 => x"0d",
          7883 => x"75",
          7884 => x"84",
          7885 => x"86",
          7886 => x"71",
          7887 => x"c0",
          7888 => x"53",
          7889 => x"38",
          7890 => x"81",
          7891 => x"51",
          7892 => x"2e",
          7893 => x"c0",
          7894 => x"55",
          7895 => x"87",
          7896 => x"08",
          7897 => x"38",
          7898 => x"87",
          7899 => x"14",
          7900 => x"82",
          7901 => x"80",
          7902 => x"38",
          7903 => x"06",
          7904 => x"38",
          7905 => x"f6",
          7906 => x"58",
          7907 => x"19",
          7908 => x"56",
          7909 => x"2e",
          7910 => x"a8",
          7911 => x"56",
          7912 => x"81",
          7913 => x"53",
          7914 => x"18",
          7915 => x"a3",
          7916 => x"e4",
          7917 => x"83",
          7918 => x"78",
          7919 => x"0c",
          7920 => x"04",
          7921 => x"18",
          7922 => x"18",
          7923 => x"19",
          7924 => x"fc",
          7925 => x"59",
          7926 => x"08",
          7927 => x"81",
          7928 => x"84",
          7929 => x"83",
          7930 => x"18",
          7931 => x"1a",
          7932 => x"1a",
          7933 => x"e4",
          7934 => x"56",
          7935 => x"27",
          7936 => x"82",
          7937 => x"74",
          7938 => x"81",
          7939 => x"38",
          7940 => x"1b",
          7941 => x"81",
          7942 => x"fc",
          7943 => x"78",
          7944 => x"75",
          7945 => x"81",
          7946 => x"38",
          7947 => x"57",
          7948 => x"09",
          7949 => x"ee",
          7950 => x"5a",
          7951 => x"56",
          7952 => x"70",
          7953 => x"34",
          7954 => x"76",
          7955 => x"d5",
          7956 => x"19",
          7957 => x"0b",
          7958 => x"34",
          7959 => x"34",
          7960 => x"b9",
          7961 => x"e1",
          7962 => x"34",
          7963 => x"bb",
          7964 => x"f2",
          7965 => x"19",
          7966 => x"0b",
          7967 => x"34",
          7968 => x"84",
          7969 => x"80",
          7970 => x"9f",
          7971 => x"18",
          7972 => x"84",
          7973 => x"74",
          7974 => x"7a",
          7975 => x"34",
          7976 => x"56",
          7977 => x"19",
          7978 => x"2a",
          7979 => x"a3",
          7980 => x"18",
          7981 => x"84",
          7982 => x"7a",
          7983 => x"74",
          7984 => x"34",
          7985 => x"56",
          7986 => x"19",
          7987 => x"2a",
          7988 => x"a7",
          7989 => x"18",
          7990 => x"70",
          7991 => x"5b",
          7992 => x"53",
          7993 => x"18",
          7994 => x"e8",
          7995 => x"19",
          7996 => x"80",
          7997 => x"33",
          7998 => x"3f",
          7999 => x"08",
          8000 => x"b7",
          8001 => x"39",
          8002 => x"60",
          8003 => x"59",
          8004 => x"76",
          8005 => x"9c",
          8006 => x"26",
          8007 => x"58",
          8008 => x"e4",
          8009 => x"0d",
          8010 => x"33",
          8011 => x"82",
          8012 => x"38",
          8013 => x"82",
          8014 => x"81",
          8015 => x"06",
          8016 => x"81",
          8017 => x"89",
          8018 => x"08",
          8019 => x"80",
          8020 => x"08",
          8021 => x"38",
          8022 => x"5c",
          8023 => x"09",
          8024 => x"de",
          8025 => x"78",
          8026 => x"52",
          8027 => x"51",
          8028 => x"84",
          8029 => x"80",
          8030 => x"ff",
          8031 => x"78",
          8032 => x"7a",
          8033 => x"79",
          8034 => x"17",
          8035 => x"81",
          8036 => x"2a",
          8037 => x"05",
          8038 => x"59",
          8039 => x"79",
          8040 => x"80",
          8041 => x"33",
          8042 => x"5d",
          8043 => x"09",
          8044 => x"b5",
          8045 => x"78",
          8046 => x"52",
          8047 => x"51",
          8048 => x"84",
          8049 => x"80",
          8050 => x"ff",
          8051 => x"78",
          8052 => x"79",
          8053 => x"7a",
          8054 => x"17",
          8055 => x"70",
          8056 => x"07",
          8057 => x"71",
          8058 => x"5d",
          8059 => x"79",
          8060 => x"76",
          8061 => x"84",
          8062 => x"8f",
          8063 => x"75",
          8064 => x"18",
          8065 => x"b4",
          8066 => x"2e",
          8067 => x"0b",
          8068 => x"71",
          8069 => x"7b",
          8070 => x"81",
          8071 => x"38",
          8072 => x"53",
          8073 => x"81",
          8074 => x"f7",
          8075 => x"b8",
          8076 => x"2e",
          8077 => x"59",
          8078 => x"b4",
          8079 => x"fd",
          8080 => x"10",
          8081 => x"77",
          8082 => x"81",
          8083 => x"33",
          8084 => x"07",
          8085 => x"0c",
          8086 => x"3d",
          8087 => x"83",
          8088 => x"06",
          8089 => x"75",
          8090 => x"18",
          8091 => x"b4",
          8092 => x"2e",
          8093 => x"0b",
          8094 => x"71",
          8095 => x"7c",
          8096 => x"81",
          8097 => x"38",
          8098 => x"53",
          8099 => x"81",
          8100 => x"f6",
          8101 => x"b8",
          8102 => x"2e",
          8103 => x"59",
          8104 => x"b4",
          8105 => x"fc",
          8106 => x"82",
          8107 => x"06",
          8108 => x"05",
          8109 => x"82",
          8110 => x"90",
          8111 => x"2b",
          8112 => x"33",
          8113 => x"88",
          8114 => x"71",
          8115 => x"fe",
          8116 => x"84",
          8117 => x"41",
          8118 => x"5a",
          8119 => x"0d",
          8120 => x"b4",
          8121 => x"b8",
          8122 => x"81",
          8123 => x"5c",
          8124 => x"81",
          8125 => x"e4",
          8126 => x"09",
          8127 => x"be",
          8128 => x"e4",
          8129 => x"34",
          8130 => x"a8",
          8131 => x"84",
          8132 => x"5b",
          8133 => x"18",
          8134 => x"84",
          8135 => x"33",
          8136 => x"2e",
          8137 => x"fd",
          8138 => x"54",
          8139 => x"a0",
          8140 => x"53",
          8141 => x"17",
          8142 => x"98",
          8143 => x"fd",
          8144 => x"54",
          8145 => x"53",
          8146 => x"53",
          8147 => x"52",
          8148 => x"3f",
          8149 => x"08",
          8150 => x"81",
          8151 => x"38",
          8152 => x"08",
          8153 => x"b4",
          8154 => x"18",
          8155 => x"7c",
          8156 => x"27",
          8157 => x"17",
          8158 => x"82",
          8159 => x"38",
          8160 => x"08",
          8161 => x"39",
          8162 => x"17",
          8163 => x"17",
          8164 => x"18",
          8165 => x"f5",
          8166 => x"5a",
          8167 => x"08",
          8168 => x"81",
          8169 => x"38",
          8170 => x"08",
          8171 => x"b4",
          8172 => x"18",
          8173 => x"b8",
          8174 => x"5e",
          8175 => x"08",
          8176 => x"38",
          8177 => x"55",
          8178 => x"09",
          8179 => x"b8",
          8180 => x"b4",
          8181 => x"18",
          8182 => x"7b",
          8183 => x"33",
          8184 => x"3f",
          8185 => x"a0",
          8186 => x"b4",
          8187 => x"b8",
          8188 => x"81",
          8189 => x"5e",
          8190 => x"81",
          8191 => x"e4",
          8192 => x"09",
          8193 => x"cb",
          8194 => x"e4",
          8195 => x"34",
          8196 => x"a8",
          8197 => x"84",
          8198 => x"5b",
          8199 => x"18",
          8200 => x"91",
          8201 => x"33",
          8202 => x"2e",
          8203 => x"fb",
          8204 => x"54",
          8205 => x"a0",
          8206 => x"53",
          8207 => x"17",
          8208 => x"90",
          8209 => x"fa",
          8210 => x"54",
          8211 => x"a0",
          8212 => x"53",
          8213 => x"17",
          8214 => x"f8",
          8215 => x"39",
          8216 => x"f9",
          8217 => x"9f",
          8218 => x"0d",
          8219 => x"5d",
          8220 => x"58",
          8221 => x"9c",
          8222 => x"1a",
          8223 => x"38",
          8224 => x"74",
          8225 => x"38",
          8226 => x"81",
          8227 => x"81",
          8228 => x"38",
          8229 => x"e4",
          8230 => x"0d",
          8231 => x"2a",
          8232 => x"05",
          8233 => x"b4",
          8234 => x"5c",
          8235 => x"86",
          8236 => x"19",
          8237 => x"5d",
          8238 => x"09",
          8239 => x"fa",
          8240 => x"77",
          8241 => x"52",
          8242 => x"51",
          8243 => x"84",
          8244 => x"80",
          8245 => x"ff",
          8246 => x"77",
          8247 => x"79",
          8248 => x"b0",
          8249 => x"83",
          8250 => x"05",
          8251 => x"ff",
          8252 => x"76",
          8253 => x"76",
          8254 => x"79",
          8255 => x"81",
          8256 => x"34",
          8257 => x"e4",
          8258 => x"0d",
          8259 => x"2e",
          8260 => x"fe",
          8261 => x"87",
          8262 => x"08",
          8263 => x"0b",
          8264 => x"58",
          8265 => x"2e",
          8266 => x"83",
          8267 => x"5b",
          8268 => x"2e",
          8269 => x"84",
          8270 => x"54",
          8271 => x"19",
          8272 => x"33",
          8273 => x"3f",
          8274 => x"08",
          8275 => x"38",
          8276 => x"5a",
          8277 => x"0c",
          8278 => x"fe",
          8279 => x"82",
          8280 => x"06",
          8281 => x"11",
          8282 => x"70",
          8283 => x"0a",
          8284 => x"0a",
          8285 => x"57",
          8286 => x"7d",
          8287 => x"2a",
          8288 => x"1d",
          8289 => x"2a",
          8290 => x"1d",
          8291 => x"2a",
          8292 => x"1d",
          8293 => x"83",
          8294 => x"e8",
          8295 => x"2a",
          8296 => x"2a",
          8297 => x"05",
          8298 => x"59",
          8299 => x"78",
          8300 => x"80",
          8301 => x"33",
          8302 => x"5d",
          8303 => x"09",
          8304 => x"d4",
          8305 => x"77",
          8306 => x"52",
          8307 => x"51",
          8308 => x"84",
          8309 => x"80",
          8310 => x"ff",
          8311 => x"77",
          8312 => x"7b",
          8313 => x"ac",
          8314 => x"ff",
          8315 => x"05",
          8316 => x"81",
          8317 => x"57",
          8318 => x"80",
          8319 => x"7a",
          8320 => x"f0",
          8321 => x"8f",
          8322 => x"56",
          8323 => x"34",
          8324 => x"1a",
          8325 => x"2a",
          8326 => x"05",
          8327 => x"b4",
          8328 => x"5f",
          8329 => x"83",
          8330 => x"54",
          8331 => x"19",
          8332 => x"1a",
          8333 => x"f0",
          8334 => x"58",
          8335 => x"08",
          8336 => x"81",
          8337 => x"38",
          8338 => x"08",
          8339 => x"b4",
          8340 => x"a8",
          8341 => x"a0",
          8342 => x"b8",
          8343 => x"5c",
          8344 => x"7a",
          8345 => x"82",
          8346 => x"74",
          8347 => x"e4",
          8348 => x"75",
          8349 => x"81",
          8350 => x"ee",
          8351 => x"b8",
          8352 => x"2e",
          8353 => x"56",
          8354 => x"b4",
          8355 => x"fc",
          8356 => x"83",
          8357 => x"b8",
          8358 => x"2a",
          8359 => x"8f",
          8360 => x"2a",
          8361 => x"f0",
          8362 => x"06",
          8363 => x"74",
          8364 => x"0b",
          8365 => x"fc",
          8366 => x"54",
          8367 => x"19",
          8368 => x"1a",
          8369 => x"ef",
          8370 => x"5a",
          8371 => x"08",
          8372 => x"81",
          8373 => x"38",
          8374 => x"08",
          8375 => x"b4",
          8376 => x"a8",
          8377 => x"a0",
          8378 => x"b8",
          8379 => x"59",
          8380 => x"77",
          8381 => x"38",
          8382 => x"55",
          8383 => x"09",
          8384 => x"bd",
          8385 => x"76",
          8386 => x"52",
          8387 => x"51",
          8388 => x"7b",
          8389 => x"39",
          8390 => x"53",
          8391 => x"53",
          8392 => x"52",
          8393 => x"3f",
          8394 => x"b8",
          8395 => x"2e",
          8396 => x"fd",
          8397 => x"b8",
          8398 => x"1a",
          8399 => x"08",
          8400 => x"08",
          8401 => x"08",
          8402 => x"08",
          8403 => x"5f",
          8404 => x"fc",
          8405 => x"19",
          8406 => x"82",
          8407 => x"06",
          8408 => x"81",
          8409 => x"53",
          8410 => x"19",
          8411 => x"e4",
          8412 => x"fc",
          8413 => x"54",
          8414 => x"19",
          8415 => x"1a",
          8416 => x"ed",
          8417 => x"5a",
          8418 => x"08",
          8419 => x"81",
          8420 => x"38",
          8421 => x"08",
          8422 => x"b4",
          8423 => x"a8",
          8424 => x"a0",
          8425 => x"b8",
          8426 => x"5f",
          8427 => x"7d",
          8428 => x"38",
          8429 => x"55",
          8430 => x"09",
          8431 => x"fa",
          8432 => x"7c",
          8433 => x"52",
          8434 => x"51",
          8435 => x"7b",
          8436 => x"39",
          8437 => x"1c",
          8438 => x"81",
          8439 => x"ec",
          8440 => x"58",
          8441 => x"7b",
          8442 => x"fe",
          8443 => x"7c",
          8444 => x"06",
          8445 => x"76",
          8446 => x"76",
          8447 => x"79",
          8448 => x"f9",
          8449 => x"58",
          8450 => x"7b",
          8451 => x"83",
          8452 => x"05",
          8453 => x"11",
          8454 => x"2b",
          8455 => x"7f",
          8456 => x"07",
          8457 => x"5d",
          8458 => x"34",
          8459 => x"56",
          8460 => x"34",
          8461 => x"5a",
          8462 => x"34",
          8463 => x"5b",
          8464 => x"34",
          8465 => x"f6",
          8466 => x"7e",
          8467 => x"5c",
          8468 => x"8a",
          8469 => x"08",
          8470 => x"2e",
          8471 => x"76",
          8472 => x"27",
          8473 => x"94",
          8474 => x"56",
          8475 => x"2e",
          8476 => x"76",
          8477 => x"93",
          8478 => x"81",
          8479 => x"19",
          8480 => x"89",
          8481 => x"75",
          8482 => x"b2",
          8483 => x"79",
          8484 => x"3f",
          8485 => x"08",
          8486 => x"d0",
          8487 => x"84",
          8488 => x"81",
          8489 => x"84",
          8490 => x"09",
          8491 => x"72",
          8492 => x"70",
          8493 => x"51",
          8494 => x"82",
          8495 => x"77",
          8496 => x"06",
          8497 => x"73",
          8498 => x"b8",
          8499 => x"3d",
          8500 => x"57",
          8501 => x"84",
          8502 => x"58",
          8503 => x"52",
          8504 => x"a4",
          8505 => x"74",
          8506 => x"08",
          8507 => x"84",
          8508 => x"55",
          8509 => x"08",
          8510 => x"38",
          8511 => x"84",
          8512 => x"26",
          8513 => x"57",
          8514 => x"81",
          8515 => x"19",
          8516 => x"83",
          8517 => x"75",
          8518 => x"ef",
          8519 => x"58",
          8520 => x"08",
          8521 => x"a0",
          8522 => x"e4",
          8523 => x"30",
          8524 => x"80",
          8525 => x"07",
          8526 => x"08",
          8527 => x"55",
          8528 => x"85",
          8529 => x"e4",
          8530 => x"9a",
          8531 => x"08",
          8532 => x"27",
          8533 => x"73",
          8534 => x"27",
          8535 => x"73",
          8536 => x"fe",
          8537 => x"80",
          8538 => x"38",
          8539 => x"52",
          8540 => x"f5",
          8541 => x"e4",
          8542 => x"e4",
          8543 => x"84",
          8544 => x"07",
          8545 => x"58",
          8546 => x"c4",
          8547 => x"e3",
          8548 => x"1a",
          8549 => x"08",
          8550 => x"1a",
          8551 => x"74",
          8552 => x"38",
          8553 => x"1a",
          8554 => x"33",
          8555 => x"79",
          8556 => x"75",
          8557 => x"b8",
          8558 => x"3d",
          8559 => x"0b",
          8560 => x"0c",
          8561 => x"04",
          8562 => x"08",
          8563 => x"39",
          8564 => x"ff",
          8565 => x"53",
          8566 => x"51",
          8567 => x"84",
          8568 => x"55",
          8569 => x"84",
          8570 => x"84",
          8571 => x"8c",
          8572 => x"ff",
          8573 => x"2e",
          8574 => x"81",
          8575 => x"39",
          8576 => x"7a",
          8577 => x"59",
          8578 => x"f0",
          8579 => x"80",
          8580 => x"9f",
          8581 => x"80",
          8582 => x"90",
          8583 => x"18",
          8584 => x"80",
          8585 => x"33",
          8586 => x"26",
          8587 => x"73",
          8588 => x"82",
          8589 => x"22",
          8590 => x"79",
          8591 => x"ac",
          8592 => x"19",
          8593 => x"19",
          8594 => x"08",
          8595 => x"72",
          8596 => x"38",
          8597 => x"13",
          8598 => x"73",
          8599 => x"17",
          8600 => x"19",
          8601 => x"75",
          8602 => x"0c",
          8603 => x"04",
          8604 => x"b8",
          8605 => x"3d",
          8606 => x"17",
          8607 => x"80",
          8608 => x"38",
          8609 => x"70",
          8610 => x"59",
          8611 => x"a5",
          8612 => x"08",
          8613 => x"fe",
          8614 => x"80",
          8615 => x"27",
          8616 => x"17",
          8617 => x"29",
          8618 => x"05",
          8619 => x"98",
          8620 => x"91",
          8621 => x"77",
          8622 => x"3f",
          8623 => x"08",
          8624 => x"e4",
          8625 => x"a4",
          8626 => x"84",
          8627 => x"27",
          8628 => x"9c",
          8629 => x"84",
          8630 => x"73",
          8631 => x"38",
          8632 => x"54",
          8633 => x"cd",
          8634 => x"39",
          8635 => x"b8",
          8636 => x"3d",
          8637 => x"3d",
          8638 => x"08",
          8639 => x"a0",
          8640 => x"57",
          8641 => x"7a",
          8642 => x"80",
          8643 => x"0c",
          8644 => x"55",
          8645 => x"80",
          8646 => x"79",
          8647 => x"5b",
          8648 => x"81",
          8649 => x"08",
          8650 => x"a9",
          8651 => x"2a",
          8652 => x"57",
          8653 => x"27",
          8654 => x"77",
          8655 => x"79",
          8656 => x"78",
          8657 => x"9c",
          8658 => x"56",
          8659 => x"e4",
          8660 => x"0d",
          8661 => x"18",
          8662 => x"22",
          8663 => x"89",
          8664 => x"7b",
          8665 => x"52",
          8666 => x"9c",
          8667 => x"e4",
          8668 => x"56",
          8669 => x"b8",
          8670 => x"d0",
          8671 => x"84",
          8672 => x"ff",
          8673 => x"9c",
          8674 => x"b8",
          8675 => x"82",
          8676 => x"80",
          8677 => x"38",
          8678 => x"52",
          8679 => x"a7",
          8680 => x"e4",
          8681 => x"56",
          8682 => x"08",
          8683 => x"9c",
          8684 => x"84",
          8685 => x"81",
          8686 => x"38",
          8687 => x"b8",
          8688 => x"2e",
          8689 => x"84",
          8690 => x"83",
          8691 => x"58",
          8692 => x"38",
          8693 => x"1a",
          8694 => x"59",
          8695 => x"75",
          8696 => x"38",
          8697 => x"76",
          8698 => x"1b",
          8699 => x"5e",
          8700 => x"0c",
          8701 => x"84",
          8702 => x"55",
          8703 => x"81",
          8704 => x"ff",
          8705 => x"f4",
          8706 => x"8a",
          8707 => x"75",
          8708 => x"80",
          8709 => x"75",
          8710 => x"52",
          8711 => x"51",
          8712 => x"84",
          8713 => x"80",
          8714 => x"16",
          8715 => x"7a",
          8716 => x"84",
          8717 => x"e4",
          8718 => x"0d",
          8719 => x"b4",
          8720 => x"b8",
          8721 => x"81",
          8722 => x"56",
          8723 => x"84",
          8724 => x"80",
          8725 => x"b8",
          8726 => x"1a",
          8727 => x"08",
          8728 => x"31",
          8729 => x"1a",
          8730 => x"e8",
          8731 => x"33",
          8732 => x"2e",
          8733 => x"fe",
          8734 => x"54",
          8735 => x"a0",
          8736 => x"53",
          8737 => x"19",
          8738 => x"c8",
          8739 => x"39",
          8740 => x"55",
          8741 => x"ff",
          8742 => x"76",
          8743 => x"06",
          8744 => x"94",
          8745 => x"1d",
          8746 => x"fe",
          8747 => x"80",
          8748 => x"27",
          8749 => x"8a",
          8750 => x"71",
          8751 => x"08",
          8752 => x"0c",
          8753 => x"39",
          8754 => x"b8",
          8755 => x"3d",
          8756 => x"3d",
          8757 => x"41",
          8758 => x"08",
          8759 => x"ff",
          8760 => x"08",
          8761 => x"75",
          8762 => x"d2",
          8763 => x"5f",
          8764 => x"58",
          8765 => x"76",
          8766 => x"38",
          8767 => x"78",
          8768 => x"78",
          8769 => x"06",
          8770 => x"81",
          8771 => x"b8",
          8772 => x"19",
          8773 => x"bd",
          8774 => x"e4",
          8775 => x"85",
          8776 => x"81",
          8777 => x"1a",
          8778 => x"76",
          8779 => x"9c",
          8780 => x"33",
          8781 => x"80",
          8782 => x"38",
          8783 => x"bf",
          8784 => x"ff",
          8785 => x"60",
          8786 => x"76",
          8787 => x"70",
          8788 => x"32",
          8789 => x"80",
          8790 => x"25",
          8791 => x"45",
          8792 => x"93",
          8793 => x"df",
          8794 => x"61",
          8795 => x"bf",
          8796 => x"2e",
          8797 => x"81",
          8798 => x"52",
          8799 => x"f6",
          8800 => x"e4",
          8801 => x"b8",
          8802 => x"b2",
          8803 => x"08",
          8804 => x"dc",
          8805 => x"b8",
          8806 => x"3d",
          8807 => x"54",
          8808 => x"53",
          8809 => x"19",
          8810 => x"a8",
          8811 => x"84",
          8812 => x"78",
          8813 => x"06",
          8814 => x"84",
          8815 => x"83",
          8816 => x"19",
          8817 => x"08",
          8818 => x"e4",
          8819 => x"7a",
          8820 => x"27",
          8821 => x"82",
          8822 => x"60",
          8823 => x"81",
          8824 => x"38",
          8825 => x"19",
          8826 => x"08",
          8827 => x"52",
          8828 => x"51",
          8829 => x"77",
          8830 => x"39",
          8831 => x"09",
          8832 => x"e7",
          8833 => x"2a",
          8834 => x"7a",
          8835 => x"38",
          8836 => x"77",
          8837 => x"70",
          8838 => x"7f",
          8839 => x"59",
          8840 => x"7d",
          8841 => x"81",
          8842 => x"5d",
          8843 => x"81",
          8844 => x"2e",
          8845 => x"fe",
          8846 => x"39",
          8847 => x"0b",
          8848 => x"7a",
          8849 => x"0c",
          8850 => x"04",
          8851 => x"df",
          8852 => x"33",
          8853 => x"2e",
          8854 => x"cb",
          8855 => x"08",
          8856 => x"9a",
          8857 => x"88",
          8858 => x"56",
          8859 => x"b7",
          8860 => x"70",
          8861 => x"8d",
          8862 => x"51",
          8863 => x"58",
          8864 => x"e4",
          8865 => x"05",
          8866 => x"71",
          8867 => x"2b",
          8868 => x"56",
          8869 => x"80",
          8870 => x"81",
          8871 => x"87",
          8872 => x"61",
          8873 => x"42",
          8874 => x"81",
          8875 => x"17",
          8876 => x"27",
          8877 => x"33",
          8878 => x"81",
          8879 => x"77",
          8880 => x"38",
          8881 => x"26",
          8882 => x"79",
          8883 => x"43",
          8884 => x"ff",
          8885 => x"ff",
          8886 => x"fd",
          8887 => x"83",
          8888 => x"ca",
          8889 => x"55",
          8890 => x"7c",
          8891 => x"55",
          8892 => x"81",
          8893 => x"80",
          8894 => x"70",
          8895 => x"33",
          8896 => x"70",
          8897 => x"ff",
          8898 => x"59",
          8899 => x"74",
          8900 => x"81",
          8901 => x"ac",
          8902 => x"84",
          8903 => x"94",
          8904 => x"ef",
          8905 => x"70",
          8906 => x"80",
          8907 => x"f5",
          8908 => x"b8",
          8909 => x"84",
          8910 => x"82",
          8911 => x"ff",
          8912 => x"ff",
          8913 => x"0c",
          8914 => x"98",
          8915 => x"80",
          8916 => x"08",
          8917 => x"cc",
          8918 => x"33",
          8919 => x"74",
          8920 => x"81",
          8921 => x"38",
          8922 => x"53",
          8923 => x"81",
          8924 => x"dc",
          8925 => x"b8",
          8926 => x"2e",
          8927 => x"56",
          8928 => x"b4",
          8929 => x"5a",
          8930 => x"38",
          8931 => x"70",
          8932 => x"76",
          8933 => x"99",
          8934 => x"33",
          8935 => x"81",
          8936 => x"58",
          8937 => x"34",
          8938 => x"2e",
          8939 => x"75",
          8940 => x"06",
          8941 => x"2e",
          8942 => x"74",
          8943 => x"75",
          8944 => x"e5",
          8945 => x"38",
          8946 => x"58",
          8947 => x"81",
          8948 => x"80",
          8949 => x"70",
          8950 => x"33",
          8951 => x"70",
          8952 => x"ff",
          8953 => x"5d",
          8954 => x"74",
          8955 => x"cd",
          8956 => x"33",
          8957 => x"76",
          8958 => x"0b",
          8959 => x"57",
          8960 => x"05",
          8961 => x"70",
          8962 => x"33",
          8963 => x"ff",
          8964 => x"42",
          8965 => x"2e",
          8966 => x"75",
          8967 => x"38",
          8968 => x"ff",
          8969 => x"0c",
          8970 => x"51",
          8971 => x"84",
          8972 => x"5a",
          8973 => x"08",
          8974 => x"8f",
          8975 => x"b8",
          8976 => x"3d",
          8977 => x"54",
          8978 => x"53",
          8979 => x"1b",
          8980 => x"80",
          8981 => x"84",
          8982 => x"78",
          8983 => x"06",
          8984 => x"84",
          8985 => x"83",
          8986 => x"1b",
          8987 => x"08",
          8988 => x"e4",
          8989 => x"78",
          8990 => x"27",
          8991 => x"82",
          8992 => x"79",
          8993 => x"81",
          8994 => x"38",
          8995 => x"1b",
          8996 => x"08",
          8997 => x"52",
          8998 => x"51",
          8999 => x"77",
          9000 => x"39",
          9001 => x"e4",
          9002 => x"33",
          9003 => x"81",
          9004 => x"60",
          9005 => x"76",
          9006 => x"06",
          9007 => x"2e",
          9008 => x"19",
          9009 => x"bf",
          9010 => x"1f",
          9011 => x"05",
          9012 => x"5f",
          9013 => x"af",
          9014 => x"55",
          9015 => x"52",
          9016 => x"92",
          9017 => x"e4",
          9018 => x"b8",
          9019 => x"2e",
          9020 => x"fe",
          9021 => x"80",
          9022 => x"38",
          9023 => x"ff",
          9024 => x"0c",
          9025 => x"8d",
          9026 => x"7e",
          9027 => x"81",
          9028 => x"8c",
          9029 => x"1a",
          9030 => x"33",
          9031 => x"07",
          9032 => x"76",
          9033 => x"78",
          9034 => x"06",
          9035 => x"05",
          9036 => x"77",
          9037 => x"e4",
          9038 => x"79",
          9039 => x"33",
          9040 => x"88",
          9041 => x"42",
          9042 => x"2e",
          9043 => x"79",
          9044 => x"ff",
          9045 => x"51",
          9046 => x"3f",
          9047 => x"08",
          9048 => x"05",
          9049 => x"43",
          9050 => x"56",
          9051 => x"3f",
          9052 => x"e4",
          9053 => x"81",
          9054 => x"38",
          9055 => x"18",
          9056 => x"27",
          9057 => x"78",
          9058 => x"2a",
          9059 => x"59",
          9060 => x"92",
          9061 => x"2e",
          9062 => x"10",
          9063 => x"22",
          9064 => x"fe",
          9065 => x"1d",
          9066 => x"06",
          9067 => x"ae",
          9068 => x"84",
          9069 => x"93",
          9070 => x"76",
          9071 => x"2e",
          9072 => x"81",
          9073 => x"94",
          9074 => x"0d",
          9075 => x"70",
          9076 => x"81",
          9077 => x"5a",
          9078 => x"56",
          9079 => x"38",
          9080 => x"08",
          9081 => x"57",
          9082 => x"2e",
          9083 => x"1d",
          9084 => x"70",
          9085 => x"5d",
          9086 => x"95",
          9087 => x"5b",
          9088 => x"7b",
          9089 => x"75",
          9090 => x"57",
          9091 => x"81",
          9092 => x"ff",
          9093 => x"ef",
          9094 => x"db",
          9095 => x"81",
          9096 => x"76",
          9097 => x"aa",
          9098 => x"0b",
          9099 => x"81",
          9100 => x"40",
          9101 => x"08",
          9102 => x"8b",
          9103 => x"57",
          9104 => x"81",
          9105 => x"76",
          9106 => x"58",
          9107 => x"55",
          9108 => x"85",
          9109 => x"c2",
          9110 => x"22",
          9111 => x"80",
          9112 => x"74",
          9113 => x"56",
          9114 => x"81",
          9115 => x"07",
          9116 => x"70",
          9117 => x"06",
          9118 => x"81",
          9119 => x"56",
          9120 => x"2e",
          9121 => x"84",
          9122 => x"57",
          9123 => x"77",
          9124 => x"38",
          9125 => x"74",
          9126 => x"02",
          9127 => x"cf",
          9128 => x"76",
          9129 => x"06",
          9130 => x"27",
          9131 => x"15",
          9132 => x"34",
          9133 => x"19",
          9134 => x"59",
          9135 => x"e3",
          9136 => x"59",
          9137 => x"34",
          9138 => x"56",
          9139 => x"a0",
          9140 => x"55",
          9141 => x"98",
          9142 => x"56",
          9143 => x"88",
          9144 => x"1a",
          9145 => x"57",
          9146 => x"09",
          9147 => x"38",
          9148 => x"a0",
          9149 => x"26",
          9150 => x"3d",
          9151 => x"05",
          9152 => x"33",
          9153 => x"74",
          9154 => x"76",
          9155 => x"38",
          9156 => x"8f",
          9157 => x"e4",
          9158 => x"81",
          9159 => x"e3",
          9160 => x"91",
          9161 => x"7a",
          9162 => x"82",
          9163 => x"b8",
          9164 => x"84",
          9165 => x"84",
          9166 => x"06",
          9167 => x"02",
          9168 => x"33",
          9169 => x"7d",
          9170 => x"05",
          9171 => x"33",
          9172 => x"81",
          9173 => x"5f",
          9174 => x"80",
          9175 => x"8d",
          9176 => x"51",
          9177 => x"3f",
          9178 => x"08",
          9179 => x"52",
          9180 => x"8c",
          9181 => x"e4",
          9182 => x"b8",
          9183 => x"82",
          9184 => x"e4",
          9185 => x"5e",
          9186 => x"08",
          9187 => x"b4",
          9188 => x"2e",
          9189 => x"83",
          9190 => x"7f",
          9191 => x"81",
          9192 => x"38",
          9193 => x"53",
          9194 => x"81",
          9195 => x"d4",
          9196 => x"b8",
          9197 => x"2e",
          9198 => x"56",
          9199 => x"b4",
          9200 => x"56",
          9201 => x"9c",
          9202 => x"33",
          9203 => x"81",
          9204 => x"c9",
          9205 => x"70",
          9206 => x"07",
          9207 => x"80",
          9208 => x"38",
          9209 => x"78",
          9210 => x"89",
          9211 => x"7d",
          9212 => x"3f",
          9213 => x"08",
          9214 => x"e4",
          9215 => x"ff",
          9216 => x"58",
          9217 => x"81",
          9218 => x"58",
          9219 => x"38",
          9220 => x"7f",
          9221 => x"98",
          9222 => x"b4",
          9223 => x"2e",
          9224 => x"1c",
          9225 => x"40",
          9226 => x"38",
          9227 => x"53",
          9228 => x"81",
          9229 => x"d3",
          9230 => x"b8",
          9231 => x"2e",
          9232 => x"57",
          9233 => x"b4",
          9234 => x"58",
          9235 => x"38",
          9236 => x"1f",
          9237 => x"80",
          9238 => x"05",
          9239 => x"15",
          9240 => x"38",
          9241 => x"1f",
          9242 => x"58",
          9243 => x"81",
          9244 => x"77",
          9245 => x"59",
          9246 => x"55",
          9247 => x"9c",
          9248 => x"1f",
          9249 => x"5e",
          9250 => x"1b",
          9251 => x"83",
          9252 => x"56",
          9253 => x"e4",
          9254 => x"0d",
          9255 => x"30",
          9256 => x"72",
          9257 => x"57",
          9258 => x"38",
          9259 => x"52",
          9260 => x"c2",
          9261 => x"e4",
          9262 => x"b8",
          9263 => x"2e",
          9264 => x"fe",
          9265 => x"54",
          9266 => x"53",
          9267 => x"18",
          9268 => x"80",
          9269 => x"e4",
          9270 => x"09",
          9271 => x"bf",
          9272 => x"e4",
          9273 => x"34",
          9274 => x"a8",
          9275 => x"55",
          9276 => x"08",
          9277 => x"82",
          9278 => x"60",
          9279 => x"ac",
          9280 => x"e4",
          9281 => x"9c",
          9282 => x"2b",
          9283 => x"71",
          9284 => x"7d",
          9285 => x"3f",
          9286 => x"08",
          9287 => x"e4",
          9288 => x"38",
          9289 => x"e4",
          9290 => x"8b",
          9291 => x"2a",
          9292 => x"29",
          9293 => x"81",
          9294 => x"57",
          9295 => x"81",
          9296 => x"19",
          9297 => x"76",
          9298 => x"81",
          9299 => x"1d",
          9300 => x"1e",
          9301 => x"56",
          9302 => x"77",
          9303 => x"83",
          9304 => x"7a",
          9305 => x"81",
          9306 => x"38",
          9307 => x"53",
          9308 => x"81",
          9309 => x"d0",
          9310 => x"b8",
          9311 => x"2e",
          9312 => x"57",
          9313 => x"b4",
          9314 => x"58",
          9315 => x"38",
          9316 => x"9c",
          9317 => x"81",
          9318 => x"5c",
          9319 => x"1c",
          9320 => x"8b",
          9321 => x"8c",
          9322 => x"9a",
          9323 => x"9b",
          9324 => x"8d",
          9325 => x"76",
          9326 => x"59",
          9327 => x"ff",
          9328 => x"78",
          9329 => x"22",
          9330 => x"58",
          9331 => x"e4",
          9332 => x"05",
          9333 => x"70",
          9334 => x"34",
          9335 => x"56",
          9336 => x"76",
          9337 => x"ff",
          9338 => x"18",
          9339 => x"27",
          9340 => x"83",
          9341 => x"81",
          9342 => x"10",
          9343 => x"58",
          9344 => x"2e",
          9345 => x"7c",
          9346 => x"0b",
          9347 => x"80",
          9348 => x"e9",
          9349 => x"b8",
          9350 => x"84",
          9351 => x"fc",
          9352 => x"ff",
          9353 => x"fe",
          9354 => x"eb",
          9355 => x"b4",
          9356 => x"b8",
          9357 => x"81",
          9358 => x"59",
          9359 => x"81",
          9360 => x"e4",
          9361 => x"38",
          9362 => x"08",
          9363 => x"b4",
          9364 => x"1d",
          9365 => x"b8",
          9366 => x"41",
          9367 => x"08",
          9368 => x"38",
          9369 => x"42",
          9370 => x"09",
          9371 => x"bc",
          9372 => x"b4",
          9373 => x"1d",
          9374 => x"78",
          9375 => x"33",
          9376 => x"3f",
          9377 => x"a4",
          9378 => x"1f",
          9379 => x"57",
          9380 => x"81",
          9381 => x"81",
          9382 => x"38",
          9383 => x"81",
          9384 => x"76",
          9385 => x"9f",
          9386 => x"39",
          9387 => x"07",
          9388 => x"39",
          9389 => x"1c",
          9390 => x"52",
          9391 => x"51",
          9392 => x"84",
          9393 => x"76",
          9394 => x"06",
          9395 => x"b8",
          9396 => x"1d",
          9397 => x"08",
          9398 => x"31",
          9399 => x"1d",
          9400 => x"38",
          9401 => x"5f",
          9402 => x"aa",
          9403 => x"e4",
          9404 => x"f8",
          9405 => x"1c",
          9406 => x"80",
          9407 => x"38",
          9408 => x"75",
          9409 => x"e8",
          9410 => x"59",
          9411 => x"2e",
          9412 => x"fa",
          9413 => x"54",
          9414 => x"a0",
          9415 => x"53",
          9416 => x"1c",
          9417 => x"ac",
          9418 => x"39",
          9419 => x"18",
          9420 => x"08",
          9421 => x"52",
          9422 => x"51",
          9423 => x"f8",
          9424 => x"3d",
          9425 => x"71",
          9426 => x"5c",
          9427 => x"1e",
          9428 => x"08",
          9429 => x"b5",
          9430 => x"08",
          9431 => x"d9",
          9432 => x"71",
          9433 => x"08",
          9434 => x"58",
          9435 => x"72",
          9436 => x"38",
          9437 => x"14",
          9438 => x"1b",
          9439 => x"7a",
          9440 => x"80",
          9441 => x"70",
          9442 => x"06",
          9443 => x"8f",
          9444 => x"83",
          9445 => x"1a",
          9446 => x"22",
          9447 => x"5b",
          9448 => x"7a",
          9449 => x"25",
          9450 => x"06",
          9451 => x"7c",
          9452 => x"57",
          9453 => x"18",
          9454 => x"89",
          9455 => x"58",
          9456 => x"16",
          9457 => x"18",
          9458 => x"74",
          9459 => x"38",
          9460 => x"81",
          9461 => x"89",
          9462 => x"70",
          9463 => x"25",
          9464 => x"77",
          9465 => x"38",
          9466 => x"8b",
          9467 => x"70",
          9468 => x"34",
          9469 => x"74",
          9470 => x"05",
          9471 => x"18",
          9472 => x"27",
          9473 => x"7c",
          9474 => x"55",
          9475 => x"16",
          9476 => x"33",
          9477 => x"38",
          9478 => x"38",
          9479 => x"1e",
          9480 => x"7c",
          9481 => x"56",
          9482 => x"17",
          9483 => x"08",
          9484 => x"55",
          9485 => x"38",
          9486 => x"34",
          9487 => x"53",
          9488 => x"88",
          9489 => x"1c",
          9490 => x"83",
          9491 => x"12",
          9492 => x"2b",
          9493 => x"07",
          9494 => x"70",
          9495 => x"2b",
          9496 => x"07",
          9497 => x"97",
          9498 => x"17",
          9499 => x"2b",
          9500 => x"5b",
          9501 => x"5b",
          9502 => x"1e",
          9503 => x"33",
          9504 => x"71",
          9505 => x"5d",
          9506 => x"1e",
          9507 => x"0d",
          9508 => x"55",
          9509 => x"77",
          9510 => x"81",
          9511 => x"58",
          9512 => x"b5",
          9513 => x"2b",
          9514 => x"81",
          9515 => x"84",
          9516 => x"83",
          9517 => x"55",
          9518 => x"27",
          9519 => x"76",
          9520 => x"38",
          9521 => x"54",
          9522 => x"74",
          9523 => x"82",
          9524 => x"80",
          9525 => x"08",
          9526 => x"19",
          9527 => x"22",
          9528 => x"79",
          9529 => x"fd",
          9530 => x"30",
          9531 => x"78",
          9532 => x"72",
          9533 => x"58",
          9534 => x"80",
          9535 => x"7a",
          9536 => x"05",
          9537 => x"8c",
          9538 => x"5b",
          9539 => x"73",
          9540 => x"5a",
          9541 => x"80",
          9542 => x"38",
          9543 => x"7e",
          9544 => x"89",
          9545 => x"bf",
          9546 => x"78",
          9547 => x"38",
          9548 => x"8c",
          9549 => x"5b",
          9550 => x"b4",
          9551 => x"2a",
          9552 => x"06",
          9553 => x"2e",
          9554 => x"14",
          9555 => x"ff",
          9556 => x"73",
          9557 => x"05",
          9558 => x"16",
          9559 => x"19",
          9560 => x"33",
          9561 => x"56",
          9562 => x"b7",
          9563 => x"39",
          9564 => x"53",
          9565 => x"7b",
          9566 => x"25",
          9567 => x"06",
          9568 => x"58",
          9569 => x"ef",
          9570 => x"70",
          9571 => x"57",
          9572 => x"70",
          9573 => x"53",
          9574 => x"83",
          9575 => x"74",
          9576 => x"81",
          9577 => x"80",
          9578 => x"38",
          9579 => x"88",
          9580 => x"33",
          9581 => x"3d",
          9582 => x"9f",
          9583 => x"a7",
          9584 => x"8c",
          9585 => x"80",
          9586 => x"70",
          9587 => x"33",
          9588 => x"81",
          9589 => x"7f",
          9590 => x"2e",
          9591 => x"83",
          9592 => x"27",
          9593 => x"10",
          9594 => x"76",
          9595 => x"57",
          9596 => x"ff",
          9597 => x"32",
          9598 => x"73",
          9599 => x"25",
          9600 => x"5b",
          9601 => x"90",
          9602 => x"dc",
          9603 => x"38",
          9604 => x"26",
          9605 => x"e4",
          9606 => x"e4",
          9607 => x"81",
          9608 => x"54",
          9609 => x"2e",
          9610 => x"73",
          9611 => x"38",
          9612 => x"33",
          9613 => x"06",
          9614 => x"73",
          9615 => x"81",
          9616 => x"7a",
          9617 => x"76",
          9618 => x"80",
          9619 => x"10",
          9620 => x"7d",
          9621 => x"62",
          9622 => x"05",
          9623 => x"54",
          9624 => x"2e",
          9625 => x"80",
          9626 => x"73",
          9627 => x"70",
          9628 => x"25",
          9629 => x"55",
          9630 => x"80",
          9631 => x"81",
          9632 => x"54",
          9633 => x"54",
          9634 => x"2e",
          9635 => x"80",
          9636 => x"30",
          9637 => x"77",
          9638 => x"57",
          9639 => x"72",
          9640 => x"73",
          9641 => x"94",
          9642 => x"55",
          9643 => x"fe",
          9644 => x"39",
          9645 => x"73",
          9646 => x"e7",
          9647 => x"e4",
          9648 => x"ff",
          9649 => x"fe",
          9650 => x"54",
          9651 => x"e4",
          9652 => x"0d",
          9653 => x"80",
          9654 => x"ff",
          9655 => x"7a",
          9656 => x"e3",
          9657 => x"ff",
          9658 => x"1d",
          9659 => x"7b",
          9660 => x"3f",
          9661 => x"08",
          9662 => x"0c",
          9663 => x"04",
          9664 => x"dc",
          9665 => x"70",
          9666 => x"07",
          9667 => x"56",
          9668 => x"a1",
          9669 => x"42",
          9670 => x"33",
          9671 => x"72",
          9672 => x"38",
          9673 => x"32",
          9674 => x"80",
          9675 => x"40",
          9676 => x"e1",
          9677 => x"0c",
          9678 => x"82",
          9679 => x"81",
          9680 => x"38",
          9681 => x"83",
          9682 => x"17",
          9683 => x"2e",
          9684 => x"17",
          9685 => x"05",
          9686 => x"a0",
          9687 => x"70",
          9688 => x"42",
          9689 => x"59",
          9690 => x"84",
          9691 => x"38",
          9692 => x"76",
          9693 => x"59",
          9694 => x"80",
          9695 => x"80",
          9696 => x"38",
          9697 => x"70",
          9698 => x"06",
          9699 => x"55",
          9700 => x"2e",
          9701 => x"73",
          9702 => x"06",
          9703 => x"2e",
          9704 => x"76",
          9705 => x"38",
          9706 => x"05",
          9707 => x"54",
          9708 => x"9d",
          9709 => x"18",
          9710 => x"ff",
          9711 => x"80",
          9712 => x"fe",
          9713 => x"5e",
          9714 => x"2e",
          9715 => x"eb",
          9716 => x"a0",
          9717 => x"a0",
          9718 => x"05",
          9719 => x"13",
          9720 => x"38",
          9721 => x"5e",
          9722 => x"70",
          9723 => x"59",
          9724 => x"74",
          9725 => x"ed",
          9726 => x"2e",
          9727 => x"74",
          9728 => x"30",
          9729 => x"55",
          9730 => x"77",
          9731 => x"38",
          9732 => x"38",
          9733 => x"7b",
          9734 => x"81",
          9735 => x"32",
          9736 => x"72",
          9737 => x"70",
          9738 => x"51",
          9739 => x"80",
          9740 => x"38",
          9741 => x"86",
          9742 => x"77",
          9743 => x"79",
          9744 => x"75",
          9745 => x"38",
          9746 => x"5b",
          9747 => x"2b",
          9748 => x"77",
          9749 => x"5d",
          9750 => x"22",
          9751 => x"56",
          9752 => x"95",
          9753 => x"33",
          9754 => x"e5",
          9755 => x"38",
          9756 => x"82",
          9757 => x"8c",
          9758 => x"8c",
          9759 => x"38",
          9760 => x"55",
          9761 => x"82",
          9762 => x"81",
          9763 => x"56",
          9764 => x"7d",
          9765 => x"7c",
          9766 => x"38",
          9767 => x"5a",
          9768 => x"81",
          9769 => x"80",
          9770 => x"79",
          9771 => x"79",
          9772 => x"7b",
          9773 => x"3f",
          9774 => x"08",
          9775 => x"56",
          9776 => x"e4",
          9777 => x"81",
          9778 => x"b8",
          9779 => x"2e",
          9780 => x"fb",
          9781 => x"85",
          9782 => x"5a",
          9783 => x"84",
          9784 => x"82",
          9785 => x"59",
          9786 => x"38",
          9787 => x"55",
          9788 => x"8c",
          9789 => x"80",
          9790 => x"39",
          9791 => x"11",
          9792 => x"22",
          9793 => x"56",
          9794 => x"f0",
          9795 => x"2e",
          9796 => x"79",
          9797 => x"fd",
          9798 => x"18",
          9799 => x"ae",
          9800 => x"06",
          9801 => x"77",
          9802 => x"ae",
          9803 => x"06",
          9804 => x"76",
          9805 => x"80",
          9806 => x"0b",
          9807 => x"53",
          9808 => x"73",
          9809 => x"a0",
          9810 => x"70",
          9811 => x"34",
          9812 => x"8a",
          9813 => x"38",
          9814 => x"58",
          9815 => x"34",
          9816 => x"bf",
          9817 => x"e4",
          9818 => x"33",
          9819 => x"b8",
          9820 => x"d6",
          9821 => x"2a",
          9822 => x"77",
          9823 => x"86",
          9824 => x"84",
          9825 => x"56",
          9826 => x"2e",
          9827 => x"90",
          9828 => x"ff",
          9829 => x"80",
          9830 => x"80",
          9831 => x"71",
          9832 => x"62",
          9833 => x"54",
          9834 => x"2e",
          9835 => x"74",
          9836 => x"7b",
          9837 => x"56",
          9838 => x"77",
          9839 => x"ae",
          9840 => x"38",
          9841 => x"76",
          9842 => x"fb",
          9843 => x"83",
          9844 => x"56",
          9845 => x"39",
          9846 => x"81",
          9847 => x"8c",
          9848 => x"77",
          9849 => x"81",
          9850 => x"38",
          9851 => x"5a",
          9852 => x"85",
          9853 => x"34",
          9854 => x"09",
          9855 => x"f6",
          9856 => x"ff",
          9857 => x"1d",
          9858 => x"84",
          9859 => x"93",
          9860 => x"74",
          9861 => x"9d",
          9862 => x"75",
          9863 => x"38",
          9864 => x"78",
          9865 => x"f7",
          9866 => x"07",
          9867 => x"57",
          9868 => x"a4",
          9869 => x"07",
          9870 => x"52",
          9871 => x"85",
          9872 => x"b8",
          9873 => x"ff",
          9874 => x"87",
          9875 => x"5a",
          9876 => x"2e",
          9877 => x"80",
          9878 => x"e4",
          9879 => x"56",
          9880 => x"ff",
          9881 => x"38",
          9882 => x"81",
          9883 => x"e4",
          9884 => x"e4",
          9885 => x"81",
          9886 => x"54",
          9887 => x"2e",
          9888 => x"73",
          9889 => x"38",
          9890 => x"33",
          9891 => x"06",
          9892 => x"73",
          9893 => x"81",
          9894 => x"78",
          9895 => x"ff",
          9896 => x"73",
          9897 => x"38",
          9898 => x"70",
          9899 => x"5f",
          9900 => x"15",
          9901 => x"26",
          9902 => x"81",
          9903 => x"ff",
          9904 => x"70",
          9905 => x"06",
          9906 => x"53",
          9907 => x"05",
          9908 => x"34",
          9909 => x"75",
          9910 => x"fc",
          9911 => x"fa",
          9912 => x"e4",
          9913 => x"81",
          9914 => x"53",
          9915 => x"ff",
          9916 => x"df",
          9917 => x"7d",
          9918 => x"5b",
          9919 => x"79",
          9920 => x"5b",
          9921 => x"cd",
          9922 => x"cc",
          9923 => x"98",
          9924 => x"2b",
          9925 => x"88",
          9926 => x"57",
          9927 => x"7b",
          9928 => x"75",
          9929 => x"54",
          9930 => x"81",
          9931 => x"a0",
          9932 => x"74",
          9933 => x"1b",
          9934 => x"39",
          9935 => x"a0",
          9936 => x"5a",
          9937 => x"2e",
          9938 => x"fa",
          9939 => x"a3",
          9940 => x"2a",
          9941 => x"7b",
          9942 => x"85",
          9943 => x"e4",
          9944 => x"0d",
          9945 => x"0d",
          9946 => x"88",
          9947 => x"05",
          9948 => x"5e",
          9949 => x"ff",
          9950 => x"59",
          9951 => x"80",
          9952 => x"38",
          9953 => x"05",
          9954 => x"9f",
          9955 => x"75",
          9956 => x"d0",
          9957 => x"38",
          9958 => x"85",
          9959 => x"d0",
          9960 => x"80",
          9961 => x"b2",
          9962 => x"10",
          9963 => x"05",
          9964 => x"5a",
          9965 => x"80",
          9966 => x"38",
          9967 => x"7f",
          9968 => x"77",
          9969 => x"7b",
          9970 => x"38",
          9971 => x"51",
          9972 => x"3f",
          9973 => x"08",
          9974 => x"70",
          9975 => x"58",
          9976 => x"86",
          9977 => x"77",
          9978 => x"5d",
          9979 => x"1d",
          9980 => x"34",
          9981 => x"17",
          9982 => x"bb",
          9983 => x"b8",
          9984 => x"ff",
          9985 => x"06",
          9986 => x"58",
          9987 => x"38",
          9988 => x"8d",
          9989 => x"2a",
          9990 => x"8a",
          9991 => x"b1",
          9992 => x"7a",
          9993 => x"ff",
          9994 => x"0c",
          9995 => x"55",
          9996 => x"53",
          9997 => x"53",
          9998 => x"52",
          9999 => x"95",
         10000 => x"e4",
         10001 => x"85",
         10002 => x"81",
         10003 => x"18",
         10004 => x"78",
         10005 => x"b7",
         10006 => x"b6",
         10007 => x"88",
         10008 => x"56",
         10009 => x"82",
         10010 => x"85",
         10011 => x"81",
         10012 => x"84",
         10013 => x"33",
         10014 => x"bf",
         10015 => x"75",
         10016 => x"cd",
         10017 => x"75",
         10018 => x"c5",
         10019 => x"17",
         10020 => x"18",
         10021 => x"2b",
         10022 => x"7c",
         10023 => x"09",
         10024 => x"ad",
         10025 => x"17",
         10026 => x"18",
         10027 => x"2b",
         10028 => x"75",
         10029 => x"dc",
         10030 => x"33",
         10031 => x"71",
         10032 => x"88",
         10033 => x"14",
         10034 => x"07",
         10035 => x"33",
         10036 => x"5a",
         10037 => x"5f",
         10038 => x"18",
         10039 => x"17",
         10040 => x"34",
         10041 => x"33",
         10042 => x"81",
         10043 => x"40",
         10044 => x"7c",
         10045 => x"d9",
         10046 => x"ff",
         10047 => x"29",
         10048 => x"33",
         10049 => x"77",
         10050 => x"77",
         10051 => x"2e",
         10052 => x"ff",
         10053 => x"42",
         10054 => x"38",
         10055 => x"33",
         10056 => x"33",
         10057 => x"07",
         10058 => x"88",
         10059 => x"75",
         10060 => x"5a",
         10061 => x"82",
         10062 => x"cc",
         10063 => x"cb",
         10064 => x"88",
         10065 => x"5c",
         10066 => x"80",
         10067 => x"11",
         10068 => x"33",
         10069 => x"71",
         10070 => x"81",
         10071 => x"72",
         10072 => x"75",
         10073 => x"53",
         10074 => x"42",
         10075 => x"c7",
         10076 => x"c6",
         10077 => x"88",
         10078 => x"58",
         10079 => x"80",
         10080 => x"38",
         10081 => x"84",
         10082 => x"79",
         10083 => x"c1",
         10084 => x"74",
         10085 => x"fd",
         10086 => x"84",
         10087 => x"56",
         10088 => x"08",
         10089 => x"a9",
         10090 => x"e4",
         10091 => x"ff",
         10092 => x"83",
         10093 => x"75",
         10094 => x"26",
         10095 => x"5d",
         10096 => x"26",
         10097 => x"81",
         10098 => x"70",
         10099 => x"7b",
         10100 => x"7b",
         10101 => x"1a",
         10102 => x"b0",
         10103 => x"59",
         10104 => x"8a",
         10105 => x"17",
         10106 => x"58",
         10107 => x"80",
         10108 => x"16",
         10109 => x"78",
         10110 => x"82",
         10111 => x"78",
         10112 => x"81",
         10113 => x"06",
         10114 => x"83",
         10115 => x"2a",
         10116 => x"78",
         10117 => x"26",
         10118 => x"0b",
         10119 => x"ff",
         10120 => x"0c",
         10121 => x"84",
         10122 => x"83",
         10123 => x"38",
         10124 => x"84",
         10125 => x"81",
         10126 => x"84",
         10127 => x"7c",
         10128 => x"84",
         10129 => x"8c",
         10130 => x"0b",
         10131 => x"80",
         10132 => x"b8",
         10133 => x"3d",
         10134 => x"0b",
         10135 => x"0c",
         10136 => x"04",
         10137 => x"11",
         10138 => x"06",
         10139 => x"74",
         10140 => x"38",
         10141 => x"81",
         10142 => x"05",
         10143 => x"7a",
         10144 => x"38",
         10145 => x"83",
         10146 => x"40",
         10147 => x"7f",
         10148 => x"70",
         10149 => x"33",
         10150 => x"05",
         10151 => x"9f",
         10152 => x"56",
         10153 => x"89",
         10154 => x"70",
         10155 => x"57",
         10156 => x"17",
         10157 => x"26",
         10158 => x"17",
         10159 => x"06",
         10160 => x"30",
         10161 => x"59",
         10162 => x"2e",
         10163 => x"85",
         10164 => x"be",
         10165 => x"32",
         10166 => x"72",
         10167 => x"7a",
         10168 => x"55",
         10169 => x"87",
         10170 => x"1c",
         10171 => x"5c",
         10172 => x"ff",
         10173 => x"56",
         10174 => x"78",
         10175 => x"cf",
         10176 => x"2a",
         10177 => x"8a",
         10178 => x"c5",
         10179 => x"fe",
         10180 => x"78",
         10181 => x"75",
         10182 => x"09",
         10183 => x"38",
         10184 => x"81",
         10185 => x"30",
         10186 => x"7b",
         10187 => x"5c",
         10188 => x"38",
         10189 => x"2e",
         10190 => x"93",
         10191 => x"5a",
         10192 => x"fa",
         10193 => x"59",
         10194 => x"2e",
         10195 => x"81",
         10196 => x"80",
         10197 => x"90",
         10198 => x"2b",
         10199 => x"19",
         10200 => x"07",
         10201 => x"fe",
         10202 => x"07",
         10203 => x"40",
         10204 => x"7a",
         10205 => x"5c",
         10206 => x"90",
         10207 => x"78",
         10208 => x"be",
         10209 => x"d9",
         10210 => x"30",
         10211 => x"72",
         10212 => x"3d",
         10213 => x"05",
         10214 => x"b6",
         10215 => x"52",
         10216 => x"78",
         10217 => x"56",
         10218 => x"80",
         10219 => x"0b",
         10220 => x"ff",
         10221 => x"0c",
         10222 => x"56",
         10223 => x"a5",
         10224 => x"7a",
         10225 => x"52",
         10226 => x"51",
         10227 => x"3f",
         10228 => x"08",
         10229 => x"38",
         10230 => x"56",
         10231 => x"0c",
         10232 => x"bf",
         10233 => x"33",
         10234 => x"88",
         10235 => x"5e",
         10236 => x"82",
         10237 => x"09",
         10238 => x"38",
         10239 => x"18",
         10240 => x"75",
         10241 => x"82",
         10242 => x"81",
         10243 => x"30",
         10244 => x"7a",
         10245 => x"42",
         10246 => x"75",
         10247 => x"b6",
         10248 => x"77",
         10249 => x"56",
         10250 => x"b8",
         10251 => x"5d",
         10252 => x"2e",
         10253 => x"83",
         10254 => x"81",
         10255 => x"bd",
         10256 => x"2e",
         10257 => x"81",
         10258 => x"5a",
         10259 => x"27",
         10260 => x"f8",
         10261 => x"0b",
         10262 => x"83",
         10263 => x"5d",
         10264 => x"81",
         10265 => x"7e",
         10266 => x"40",
         10267 => x"31",
         10268 => x"52",
         10269 => x"80",
         10270 => x"38",
         10271 => x"e1",
         10272 => x"81",
         10273 => x"e4",
         10274 => x"58",
         10275 => x"05",
         10276 => x"70",
         10277 => x"33",
         10278 => x"ff",
         10279 => x"42",
         10280 => x"2e",
         10281 => x"75",
         10282 => x"38",
         10283 => x"f3",
         10284 => x"7c",
         10285 => x"77",
         10286 => x"0c",
         10287 => x"04",
         10288 => x"80",
         10289 => x"38",
         10290 => x"8a",
         10291 => x"98",
         10292 => x"ff",
         10293 => x"0b",
         10294 => x"0c",
         10295 => x"04",
         10296 => x"ee",
         10297 => x"94",
         10298 => x"78",
         10299 => x"5a",
         10300 => x"81",
         10301 => x"71",
         10302 => x"1b",
         10303 => x"5f",
         10304 => x"83",
         10305 => x"80",
         10306 => x"85",
         10307 => x"18",
         10308 => x"5c",
         10309 => x"70",
         10310 => x"33",
         10311 => x"05",
         10312 => x"71",
         10313 => x"5b",
         10314 => x"77",
         10315 => x"91",
         10316 => x"2e",
         10317 => x"3d",
         10318 => x"83",
         10319 => x"39",
         10320 => x"c6",
         10321 => x"17",
         10322 => x"18",
         10323 => x"2b",
         10324 => x"75",
         10325 => x"81",
         10326 => x"38",
         10327 => x"80",
         10328 => x"08",
         10329 => x"38",
         10330 => x"5b",
         10331 => x"09",
         10332 => x"9b",
         10333 => x"77",
         10334 => x"52",
         10335 => x"51",
         10336 => x"3f",
         10337 => x"08",
         10338 => x"38",
         10339 => x"5a",
         10340 => x"0c",
         10341 => x"38",
         10342 => x"34",
         10343 => x"33",
         10344 => x"33",
         10345 => x"07",
         10346 => x"82",
         10347 => x"09",
         10348 => x"fc",
         10349 => x"83",
         10350 => x"12",
         10351 => x"2b",
         10352 => x"07",
         10353 => x"70",
         10354 => x"2b",
         10355 => x"07",
         10356 => x"45",
         10357 => x"77",
         10358 => x"a4",
         10359 => x"81",
         10360 => x"38",
         10361 => x"83",
         10362 => x"12",
         10363 => x"2b",
         10364 => x"07",
         10365 => x"70",
         10366 => x"2b",
         10367 => x"07",
         10368 => x"5b",
         10369 => x"60",
         10370 => x"e4",
         10371 => x"81",
         10372 => x"38",
         10373 => x"83",
         10374 => x"12",
         10375 => x"2b",
         10376 => x"07",
         10377 => x"70",
         10378 => x"2b",
         10379 => x"07",
         10380 => x"5d",
         10381 => x"83",
         10382 => x"12",
         10383 => x"2b",
         10384 => x"07",
         10385 => x"70",
         10386 => x"2b",
         10387 => x"07",
         10388 => x"0c",
         10389 => x"46",
         10390 => x"45",
         10391 => x"7c",
         10392 => x"d0",
         10393 => x"05",
         10394 => x"d0",
         10395 => x"86",
         10396 => x"d0",
         10397 => x"18",
         10398 => x"98",
         10399 => x"cf",
         10400 => x"24",
         10401 => x"7b",
         10402 => x"56",
         10403 => x"75",
         10404 => x"08",
         10405 => x"70",
         10406 => x"33",
         10407 => x"af",
         10408 => x"b8",
         10409 => x"2e",
         10410 => x"81",
         10411 => x"b8",
         10412 => x"18",
         10413 => x"08",
         10414 => x"31",
         10415 => x"18",
         10416 => x"38",
         10417 => x"41",
         10418 => x"81",
         10419 => x"b8",
         10420 => x"fd",
         10421 => x"56",
         10422 => x"f3",
         10423 => x"0b",
         10424 => x"83",
         10425 => x"5a",
         10426 => x"39",
         10427 => x"33",
         10428 => x"33",
         10429 => x"07",
         10430 => x"58",
         10431 => x"38",
         10432 => x"42",
         10433 => x"38",
         10434 => x"83",
         10435 => x"12",
         10436 => x"2b",
         10437 => x"07",
         10438 => x"70",
         10439 => x"2b",
         10440 => x"07",
         10441 => x"5a",
         10442 => x"5a",
         10443 => x"59",
         10444 => x"39",
         10445 => x"80",
         10446 => x"38",
         10447 => x"e3",
         10448 => x"2e",
         10449 => x"93",
         10450 => x"5a",
         10451 => x"f2",
         10452 => x"79",
         10453 => x"fc",
         10454 => x"54",
         10455 => x"a0",
         10456 => x"53",
         10457 => x"17",
         10458 => x"ad",
         10459 => x"85",
         10460 => x"0d",
         10461 => x"05",
         10462 => x"43",
         10463 => x"57",
         10464 => x"5a",
         10465 => x"2e",
         10466 => x"78",
         10467 => x"5a",
         10468 => x"26",
         10469 => x"ba",
         10470 => x"38",
         10471 => x"74",
         10472 => x"d9",
         10473 => x"c0",
         10474 => x"74",
         10475 => x"38",
         10476 => x"84",
         10477 => x"70",
         10478 => x"73",
         10479 => x"38",
         10480 => x"62",
         10481 => x"2e",
         10482 => x"74",
         10483 => x"73",
         10484 => x"54",
         10485 => x"92",
         10486 => x"93",
         10487 => x"84",
         10488 => x"81",
         10489 => x"e4",
         10490 => x"84",
         10491 => x"92",
         10492 => x"8b",
         10493 => x"e4",
         10494 => x"0d",
         10495 => x"d0",
         10496 => x"ff",
         10497 => x"57",
         10498 => x"91",
         10499 => x"77",
         10500 => x"d0",
         10501 => x"77",
         10502 => x"f7",
         10503 => x"08",
         10504 => x"5e",
         10505 => x"08",
         10506 => x"79",
         10507 => x"5b",
         10508 => x"81",
         10509 => x"ff",
         10510 => x"57",
         10511 => x"26",
         10512 => x"15",
         10513 => x"06",
         10514 => x"9f",
         10515 => x"99",
         10516 => x"e0",
         10517 => x"ff",
         10518 => x"74",
         10519 => x"2a",
         10520 => x"76",
         10521 => x"06",
         10522 => x"ff",
         10523 => x"79",
         10524 => x"70",
         10525 => x"2a",
         10526 => x"57",
         10527 => x"2e",
         10528 => x"1b",
         10529 => x"5b",
         10530 => x"ff",
         10531 => x"54",
         10532 => x"7a",
         10533 => x"38",
         10534 => x"0c",
         10535 => x"39",
         10536 => x"6c",
         10537 => x"80",
         10538 => x"56",
         10539 => x"78",
         10540 => x"38",
         10541 => x"70",
         10542 => x"cc",
         10543 => x"3d",
         10544 => x"58",
         10545 => x"84",
         10546 => x"57",
         10547 => x"08",
         10548 => x"38",
         10549 => x"76",
         10550 => x"b8",
         10551 => x"3d",
         10552 => x"40",
         10553 => x"3d",
         10554 => x"e1",
         10555 => x"b8",
         10556 => x"84",
         10557 => x"80",
         10558 => x"38",
         10559 => x"5d",
         10560 => x"81",
         10561 => x"80",
         10562 => x"38",
         10563 => x"83",
         10564 => x"88",
         10565 => x"ff",
         10566 => x"83",
         10567 => x"5b",
         10568 => x"81",
         10569 => x"9b",
         10570 => x"12",
         10571 => x"2b",
         10572 => x"33",
         10573 => x"5e",
         10574 => x"2e",
         10575 => x"80",
         10576 => x"34",
         10577 => x"17",
         10578 => x"90",
         10579 => x"cc",
         10580 => x"34",
         10581 => x"0b",
         10582 => x"7e",
         10583 => x"80",
         10584 => x"34",
         10585 => x"17",
         10586 => x"5d",
         10587 => x"84",
         10588 => x"5b",
         10589 => x"1c",
         10590 => x"9d",
         10591 => x"0b",
         10592 => x"80",
         10593 => x"34",
         10594 => x"0b",
         10595 => x"7b",
         10596 => x"e2",
         10597 => x"11",
         10598 => x"08",
         10599 => x"57",
         10600 => x"89",
         10601 => x"08",
         10602 => x"8a",
         10603 => x"80",
         10604 => x"a3",
         10605 => x"e7",
         10606 => x"98",
         10607 => x"7b",
         10608 => x"b8",
         10609 => x"9c",
         10610 => x"7c",
         10611 => x"76",
         10612 => x"02",
         10613 => x"33",
         10614 => x"81",
         10615 => x"7b",
         10616 => x"77",
         10617 => x"06",
         10618 => x"2e",
         10619 => x"81",
         10620 => x"81",
         10621 => x"83",
         10622 => x"56",
         10623 => x"86",
         10624 => x"c0",
         10625 => x"b4",
         10626 => x"1b",
         10627 => x"1b",
         10628 => x"11",
         10629 => x"33",
         10630 => x"07",
         10631 => x"5e",
         10632 => x"7b",
         10633 => x"f1",
         10634 => x"1a",
         10635 => x"83",
         10636 => x"12",
         10637 => x"2b",
         10638 => x"07",
         10639 => x"70",
         10640 => x"2b",
         10641 => x"07",
         10642 => x"05",
         10643 => x"0c",
         10644 => x"59",
         10645 => x"86",
         10646 => x"1a",
         10647 => x"1a",
         10648 => x"91",
         10649 => x"0b",
         10650 => x"77",
         10651 => x"06",
         10652 => x"2e",
         10653 => x"75",
         10654 => x"f1",
         10655 => x"1a",
         10656 => x"22",
         10657 => x"7c",
         10658 => x"76",
         10659 => x"07",
         10660 => x"5b",
         10661 => x"84",
         10662 => x"70",
         10663 => x"5b",
         10664 => x"84",
         10665 => x"52",
         10666 => x"ac",
         10667 => x"b8",
         10668 => x"84",
         10669 => x"81",
         10670 => x"82",
         10671 => x"e4",
         10672 => x"80",
         10673 => x"7a",
         10674 => x"39",
         10675 => x"05",
         10676 => x"5e",
         10677 => x"77",
         10678 => x"06",
         10679 => x"2e",
         10680 => x"88",
         10681 => x"0c",
         10682 => x"87",
         10683 => x"0c",
         10684 => x"84",
         10685 => x"0c",
         10686 => x"79",
         10687 => x"3f",
         10688 => x"08",
         10689 => x"59",
         10690 => x"c8",
         10691 => x"39",
         10692 => x"31",
         10693 => x"f3",
         10694 => x"33",
         10695 => x"71",
         10696 => x"90",
         10697 => x"07",
         10698 => x"fd",
         10699 => x"55",
         10700 => x"81",
         10701 => x"52",
         10702 => x"ab",
         10703 => x"b8",
         10704 => x"84",
         10705 => x"80",
         10706 => x"38",
         10707 => x"08",
         10708 => x"d9",
         10709 => x"e4",
         10710 => x"83",
         10711 => x"53",
         10712 => x"51",
         10713 => x"3f",
         10714 => x"08",
         10715 => x"9c",
         10716 => x"11",
         10717 => x"58",
         10718 => x"75",
         10719 => x"38",
         10720 => x"18",
         10721 => x"33",
         10722 => x"74",
         10723 => x"7c",
         10724 => x"26",
         10725 => x"80",
         10726 => x"0b",
         10727 => x"80",
         10728 => x"34",
         10729 => x"95",
         10730 => x"17",
         10731 => x"2b",
         10732 => x"07",
         10733 => x"56",
         10734 => x"8e",
         10735 => x"0b",
         10736 => x"a1",
         10737 => x"34",
         10738 => x"91",
         10739 => x"56",
         10740 => x"17",
         10741 => x"57",
         10742 => x"9a",
         10743 => x"0b",
         10744 => x"7d",
         10745 => x"83",
         10746 => x"06",
         10747 => x"ff",
         10748 => x"7f",
         10749 => x"59",
         10750 => x"16",
         10751 => x"ae",
         10752 => x"33",
         10753 => x"2e",
         10754 => x"b5",
         10755 => x"7d",
         10756 => x"52",
         10757 => x"51",
         10758 => x"3f",
         10759 => x"08",
         10760 => x"38",
         10761 => x"5b",
         10762 => x"0c",
         10763 => x"ff",
         10764 => x"0c",
         10765 => x"2e",
         10766 => x"80",
         10767 => x"97",
         10768 => x"b4",
         10769 => x"b8",
         10770 => x"81",
         10771 => x"5a",
         10772 => x"3f",
         10773 => x"08",
         10774 => x"81",
         10775 => x"38",
         10776 => x"08",
         10777 => x"b4",
         10778 => x"17",
         10779 => x"b8",
         10780 => x"55",
         10781 => x"08",
         10782 => x"38",
         10783 => x"55",
         10784 => x"09",
         10785 => x"85",
         10786 => x"b4",
         10787 => x"17",
         10788 => x"79",
         10789 => x"33",
         10790 => x"b8",
         10791 => x"fe",
         10792 => x"94",
         10793 => x"56",
         10794 => x"77",
         10795 => x"76",
         10796 => x"75",
         10797 => x"5a",
         10798 => x"f8",
         10799 => x"fe",
         10800 => x"08",
         10801 => x"59",
         10802 => x"27",
         10803 => x"8a",
         10804 => x"71",
         10805 => x"08",
         10806 => x"74",
         10807 => x"cd",
         10808 => x"2a",
         10809 => x"0c",
         10810 => x"ed",
         10811 => x"1a",
         10812 => x"f7",
         10813 => x"57",
         10814 => x"f7",
         10815 => x"b8",
         10816 => x"80",
         10817 => x"cf",
         10818 => x"57",
         10819 => x"39",
         10820 => x"62",
         10821 => x"40",
         10822 => x"80",
         10823 => x"57",
         10824 => x"9f",
         10825 => x"56",
         10826 => x"97",
         10827 => x"55",
         10828 => x"8f",
         10829 => x"22",
         10830 => x"59",
         10831 => x"2e",
         10832 => x"80",
         10833 => x"76",
         10834 => x"8c",
         10835 => x"33",
         10836 => x"84",
         10837 => x"33",
         10838 => x"87",
         10839 => x"2e",
         10840 => x"94",
         10841 => x"1b",
         10842 => x"56",
         10843 => x"26",
         10844 => x"7b",
         10845 => x"d5",
         10846 => x"75",
         10847 => x"5b",
         10848 => x"38",
         10849 => x"ff",
         10850 => x"2a",
         10851 => x"9b",
         10852 => x"d3",
         10853 => x"08",
         10854 => x"27",
         10855 => x"74",
         10856 => x"f0",
         10857 => x"1b",
         10858 => x"98",
         10859 => x"05",
         10860 => x"fe",
         10861 => x"76",
         10862 => x"e7",
         10863 => x"22",
         10864 => x"b0",
         10865 => x"56",
         10866 => x"2e",
         10867 => x"7a",
         10868 => x"2a",
         10869 => x"80",
         10870 => x"38",
         10871 => x"75",
         10872 => x"38",
         10873 => x"58",
         10874 => x"53",
         10875 => x"19",
         10876 => x"9f",
         10877 => x"b8",
         10878 => x"98",
         10879 => x"11",
         10880 => x"75",
         10881 => x"38",
         10882 => x"77",
         10883 => x"78",
         10884 => x"84",
         10885 => x"29",
         10886 => x"58",
         10887 => x"70",
         10888 => x"33",
         10889 => x"05",
         10890 => x"15",
         10891 => x"38",
         10892 => x"58",
         10893 => x"7e",
         10894 => x"0c",
         10895 => x"1c",
         10896 => x"59",
         10897 => x"5e",
         10898 => x"af",
         10899 => x"75",
         10900 => x"0c",
         10901 => x"04",
         10902 => x"e4",
         10903 => x"0d",
         10904 => x"fe",
         10905 => x"1a",
         10906 => x"83",
         10907 => x"80",
         10908 => x"5b",
         10909 => x"83",
         10910 => x"76",
         10911 => x"08",
         10912 => x"38",
         10913 => x"1a",
         10914 => x"41",
         10915 => x"2e",
         10916 => x"80",
         10917 => x"54",
         10918 => x"19",
         10919 => x"33",
         10920 => x"b1",
         10921 => x"e4",
         10922 => x"85",
         10923 => x"81",
         10924 => x"1a",
         10925 => x"dc",
         10926 => x"1b",
         10927 => x"06",
         10928 => x"5a",
         10929 => x"56",
         10930 => x"2e",
         10931 => x"74",
         10932 => x"56",
         10933 => x"81",
         10934 => x"ff",
         10935 => x"80",
         10936 => x"38",
         10937 => x"05",
         10938 => x"70",
         10939 => x"34",
         10940 => x"75",
         10941 => x"bc",
         10942 => x"b4",
         10943 => x"b8",
         10944 => x"81",
         10945 => x"40",
         10946 => x"3f",
         10947 => x"b8",
         10948 => x"2e",
         10949 => x"ff",
         10950 => x"b8",
         10951 => x"1a",
         10952 => x"08",
         10953 => x"31",
         10954 => x"08",
         10955 => x"a0",
         10956 => x"fe",
         10957 => x"19",
         10958 => x"82",
         10959 => x"06",
         10960 => x"81",
         10961 => x"08",
         10962 => x"05",
         10963 => x"81",
         10964 => x"ff",
         10965 => x"7e",
         10966 => x"39",
         10967 => x"0c",
         10968 => x"56",
         10969 => x"98",
         10970 => x"79",
         10971 => x"98",
         10972 => x"e4",
         10973 => x"a1",
         10974 => x"33",
         10975 => x"83",
         10976 => x"e4",
         10977 => x"55",
         10978 => x"38",
         10979 => x"56",
         10980 => x"39",
         10981 => x"1b",
         10982 => x"84",
         10983 => x"92",
         10984 => x"82",
         10985 => x"34",
         10986 => x"b8",
         10987 => x"3d",
         10988 => x"3d",
         10989 => x"67",
         10990 => x"5c",
         10991 => x"0c",
         10992 => x"80",
         10993 => x"79",
         10994 => x"80",
         10995 => x"75",
         10996 => x"80",
         10997 => x"86",
         10998 => x"1b",
         10999 => x"78",
         11000 => x"fd",
         11001 => x"74",
         11002 => x"76",
         11003 => x"91",
         11004 => x"74",
         11005 => x"90",
         11006 => x"81",
         11007 => x"58",
         11008 => x"76",
         11009 => x"a1",
         11010 => x"08",
         11011 => x"57",
         11012 => x"84",
         11013 => x"5b",
         11014 => x"82",
         11015 => x"83",
         11016 => x"7e",
         11017 => x"60",
         11018 => x"ff",
         11019 => x"2a",
         11020 => x"78",
         11021 => x"84",
         11022 => x"1a",
         11023 => x"80",
         11024 => x"38",
         11025 => x"86",
         11026 => x"ff",
         11027 => x"38",
         11028 => x"0c",
         11029 => x"85",
         11030 => x"1b",
         11031 => x"b4",
         11032 => x"1b",
         11033 => x"d3",
         11034 => x"08",
         11035 => x"17",
         11036 => x"58",
         11037 => x"27",
         11038 => x"8a",
         11039 => x"79",
         11040 => x"08",
         11041 => x"74",
         11042 => x"de",
         11043 => x"7b",
         11044 => x"5c",
         11045 => x"83",
         11046 => x"19",
         11047 => x"27",
         11048 => x"79",
         11049 => x"54",
         11050 => x"52",
         11051 => x"51",
         11052 => x"3f",
         11053 => x"08",
         11054 => x"60",
         11055 => x"7d",
         11056 => x"74",
         11057 => x"38",
         11058 => x"b8",
         11059 => x"29",
         11060 => x"56",
         11061 => x"05",
         11062 => x"70",
         11063 => x"34",
         11064 => x"75",
         11065 => x"59",
         11066 => x"34",
         11067 => x"59",
         11068 => x"7e",
         11069 => x"0c",
         11070 => x"1c",
         11071 => x"71",
         11072 => x"8c",
         11073 => x"5a",
         11074 => x"75",
         11075 => x"38",
         11076 => x"8c",
         11077 => x"fe",
         11078 => x"1a",
         11079 => x"80",
         11080 => x"7a",
         11081 => x"80",
         11082 => x"b8",
         11083 => x"3d",
         11084 => x"84",
         11085 => x"92",
         11086 => x"83",
         11087 => x"74",
         11088 => x"60",
         11089 => x"39",
         11090 => x"08",
         11091 => x"83",
         11092 => x"80",
         11093 => x"5c",
         11094 => x"83",
         11095 => x"77",
         11096 => x"08",
         11097 => x"38",
         11098 => x"17",
         11099 => x"41",
         11100 => x"2e",
         11101 => x"80",
         11102 => x"54",
         11103 => x"16",
         11104 => x"33",
         11105 => x"cd",
         11106 => x"e4",
         11107 => x"85",
         11108 => x"81",
         11109 => x"17",
         11110 => x"bf",
         11111 => x"1b",
         11112 => x"06",
         11113 => x"b8",
         11114 => x"56",
         11115 => x"2e",
         11116 => x"70",
         11117 => x"33",
         11118 => x"05",
         11119 => x"16",
         11120 => x"38",
         11121 => x"0b",
         11122 => x"fe",
         11123 => x"54",
         11124 => x"53",
         11125 => x"53",
         11126 => x"52",
         11127 => x"f4",
         11128 => x"84",
         11129 => x"7f",
         11130 => x"06",
         11131 => x"84",
         11132 => x"83",
         11133 => x"16",
         11134 => x"08",
         11135 => x"e4",
         11136 => x"74",
         11137 => x"27",
         11138 => x"82",
         11139 => x"74",
         11140 => x"81",
         11141 => x"38",
         11142 => x"16",
         11143 => x"08",
         11144 => x"52",
         11145 => x"51",
         11146 => x"3f",
         11147 => x"ca",
         11148 => x"08",
         11149 => x"08",
         11150 => x"38",
         11151 => x"40",
         11152 => x"38",
         11153 => x"12",
         11154 => x"08",
         11155 => x"7c",
         11156 => x"58",
         11157 => x"98",
         11158 => x"79",
         11159 => x"e7",
         11160 => x"e4",
         11161 => x"b8",
         11162 => x"d8",
         11163 => x"33",
         11164 => x"39",
         11165 => x"51",
         11166 => x"3f",
         11167 => x"08",
         11168 => x"e4",
         11169 => x"38",
         11170 => x"54",
         11171 => x"53",
         11172 => x"53",
         11173 => x"52",
         11174 => x"b8",
         11175 => x"e4",
         11176 => x"38",
         11177 => x"08",
         11178 => x"b4",
         11179 => x"17",
         11180 => x"77",
         11181 => x"27",
         11182 => x"82",
         11183 => x"7b",
         11184 => x"81",
         11185 => x"38",
         11186 => x"16",
         11187 => x"08",
         11188 => x"52",
         11189 => x"51",
         11190 => x"3f",
         11191 => x"89",
         11192 => x"33",
         11193 => x"9b",
         11194 => x"e4",
         11195 => x"55",
         11196 => x"38",
         11197 => x"56",
         11198 => x"39",
         11199 => x"16",
         11200 => x"16",
         11201 => x"17",
         11202 => x"ff",
         11203 => x"84",
         11204 => x"80",
         11205 => x"b8",
         11206 => x"17",
         11207 => x"08",
         11208 => x"31",
         11209 => x"17",
         11210 => x"98",
         11211 => x"33",
         11212 => x"2e",
         11213 => x"fe",
         11214 => x"54",
         11215 => x"a0",
         11216 => x"53",
         11217 => x"16",
         11218 => x"96",
         11219 => x"7c",
         11220 => x"94",
         11221 => x"56",
         11222 => x"81",
         11223 => x"34",
         11224 => x"b8",
         11225 => x"3d",
         11226 => x"0b",
         11227 => x"82",
         11228 => x"e4",
         11229 => x"0d",
         11230 => x"0d",
         11231 => x"5a",
         11232 => x"9f",
         11233 => x"56",
         11234 => x"97",
         11235 => x"55",
         11236 => x"8f",
         11237 => x"22",
         11238 => x"58",
         11239 => x"2e",
         11240 => x"80",
         11241 => x"79",
         11242 => x"d8",
         11243 => x"33",
         11244 => x"81",
         11245 => x"7a",
         11246 => x"c8",
         11247 => x"19",
         11248 => x"b4",
         11249 => x"2e",
         11250 => x"17",
         11251 => x"81",
         11252 => x"54",
         11253 => x"17",
         11254 => x"33",
         11255 => x"f5",
         11256 => x"e4",
         11257 => x"85",
         11258 => x"81",
         11259 => x"18",
         11260 => x"90",
         11261 => x"08",
         11262 => x"a0",
         11263 => x"78",
         11264 => x"77",
         11265 => x"08",
         11266 => x"ff",
         11267 => x"56",
         11268 => x"34",
         11269 => x"5a",
         11270 => x"34",
         11271 => x"33",
         11272 => x"56",
         11273 => x"2e",
         11274 => x"8c",
         11275 => x"74",
         11276 => x"88",
         11277 => x"9d",
         11278 => x"90",
         11279 => x"9e",
         11280 => x"98",
         11281 => x"9f",
         11282 => x"7a",
         11283 => x"97",
         11284 => x"0b",
         11285 => x"80",
         11286 => x"18",
         11287 => x"92",
         11288 => x"0b",
         11289 => x"7b",
         11290 => x"83",
         11291 => x"51",
         11292 => x"3f",
         11293 => x"08",
         11294 => x"81",
         11295 => x"56",
         11296 => x"34",
         11297 => x"e4",
         11298 => x"0d",
         11299 => x"b4",
         11300 => x"b8",
         11301 => x"81",
         11302 => x"5b",
         11303 => x"3f",
         11304 => x"b8",
         11305 => x"c9",
         11306 => x"e4",
         11307 => x"34",
         11308 => x"a8",
         11309 => x"84",
         11310 => x"57",
         11311 => x"18",
         11312 => x"8e",
         11313 => x"33",
         11314 => x"2e",
         11315 => x"fe",
         11316 => x"54",
         11317 => x"a0",
         11318 => x"53",
         11319 => x"17",
         11320 => x"92",
         11321 => x"56",
         11322 => x"78",
         11323 => x"74",
         11324 => x"74",
         11325 => x"75",
         11326 => x"8c",
         11327 => x"74",
         11328 => x"88",
         11329 => x"9d",
         11330 => x"90",
         11331 => x"9e",
         11332 => x"98",
         11333 => x"9f",
         11334 => x"7a",
         11335 => x"97",
         11336 => x"0b",
         11337 => x"80",
         11338 => x"18",
         11339 => x"92",
         11340 => x"0b",
         11341 => x"7b",
         11342 => x"83",
         11343 => x"51",
         11344 => x"3f",
         11345 => x"08",
         11346 => x"81",
         11347 => x"56",
         11348 => x"34",
         11349 => x"81",
         11350 => x"ff",
         11351 => x"84",
         11352 => x"81",
         11353 => x"fc",
         11354 => x"78",
         11355 => x"fc",
         11356 => x"3d",
         11357 => x"52",
         11358 => x"3f",
         11359 => x"08",
         11360 => x"e4",
         11361 => x"89",
         11362 => x"2e",
         11363 => x"08",
         11364 => x"2e",
         11365 => x"33",
         11366 => x"2e",
         11367 => x"13",
         11368 => x"22",
         11369 => x"77",
         11370 => x"80",
         11371 => x"75",
         11372 => x"38",
         11373 => x"73",
         11374 => x"0c",
         11375 => x"04",
         11376 => x"51",
         11377 => x"3f",
         11378 => x"08",
         11379 => x"72",
         11380 => x"75",
         11381 => x"d5",
         11382 => x"0d",
         11383 => x"5b",
         11384 => x"80",
         11385 => x"75",
         11386 => x"57",
         11387 => x"26",
         11388 => x"ba",
         11389 => x"70",
         11390 => x"ba",
         11391 => x"84",
         11392 => x"51",
         11393 => x"90",
         11394 => x"d0",
         11395 => x"0b",
         11396 => x"0c",
         11397 => x"04",
         11398 => x"b8",
         11399 => x"3d",
         11400 => x"33",
         11401 => x"81",
         11402 => x"53",
         11403 => x"26",
         11404 => x"19",
         11405 => x"06",
         11406 => x"54",
         11407 => x"80",
         11408 => x"0b",
         11409 => x"5b",
         11410 => x"79",
         11411 => x"70",
         11412 => x"33",
         11413 => x"05",
         11414 => x"9f",
         11415 => x"52",
         11416 => x"89",
         11417 => x"70",
         11418 => x"53",
         11419 => x"13",
         11420 => x"26",
         11421 => x"13",
         11422 => x"06",
         11423 => x"30",
         11424 => x"55",
         11425 => x"2e",
         11426 => x"85",
         11427 => x"be",
         11428 => x"32",
         11429 => x"72",
         11430 => x"76",
         11431 => x"52",
         11432 => x"92",
         11433 => x"84",
         11434 => x"83",
         11435 => x"99",
         11436 => x"fe",
         11437 => x"83",
         11438 => x"77",
         11439 => x"fe",
         11440 => x"3d",
         11441 => x"98",
         11442 => x"52",
         11443 => x"d1",
         11444 => x"b8",
         11445 => x"84",
         11446 => x"80",
         11447 => x"74",
         11448 => x"0c",
         11449 => x"04",
         11450 => x"52",
         11451 => x"05",
         11452 => x"3f",
         11453 => x"08",
         11454 => x"e4",
         11455 => x"38",
         11456 => x"05",
         11457 => x"2b",
         11458 => x"77",
         11459 => x"38",
         11460 => x"33",
         11461 => x"81",
         11462 => x"75",
         11463 => x"38",
         11464 => x"11",
         11465 => x"33",
         11466 => x"07",
         11467 => x"5a",
         11468 => x"79",
         11469 => x"38",
         11470 => x"0c",
         11471 => x"e4",
         11472 => x"0d",
         11473 => x"e4",
         11474 => x"09",
         11475 => x"8f",
         11476 => x"84",
         11477 => x"98",
         11478 => x"95",
         11479 => x"17",
         11480 => x"2b",
         11481 => x"07",
         11482 => x"1b",
         11483 => x"cc",
         11484 => x"98",
         11485 => x"74",
         11486 => x"0c",
         11487 => x"04",
         11488 => x"0d",
         11489 => x"08",
         11490 => x"08",
         11491 => x"7c",
         11492 => x"80",
         11493 => x"b4",
         11494 => x"e5",
         11495 => x"c5",
         11496 => x"e4",
         11497 => x"b8",
         11498 => x"c8",
         11499 => x"d9",
         11500 => x"61",
         11501 => x"80",
         11502 => x"58",
         11503 => x"08",
         11504 => x"80",
         11505 => x"38",
         11506 => x"98",
         11507 => x"a0",
         11508 => x"ff",
         11509 => x"84",
         11510 => x"59",
         11511 => x"08",
         11512 => x"60",
         11513 => x"08",
         11514 => x"16",
         11515 => x"b1",
         11516 => x"e4",
         11517 => x"33",
         11518 => x"83",
         11519 => x"54",
         11520 => x"16",
         11521 => x"33",
         11522 => x"c9",
         11523 => x"e4",
         11524 => x"85",
         11525 => x"81",
         11526 => x"17",
         11527 => x"d4",
         11528 => x"3d",
         11529 => x"33",
         11530 => x"71",
         11531 => x"63",
         11532 => x"40",
         11533 => x"78",
         11534 => x"da",
         11535 => x"db",
         11536 => x"52",
         11537 => x"a3",
         11538 => x"b8",
         11539 => x"84",
         11540 => x"82",
         11541 => x"52",
         11542 => x"a8",
         11543 => x"b8",
         11544 => x"84",
         11545 => x"bb",
         11546 => x"3d",
         11547 => x"33",
         11548 => x"71",
         11549 => x"63",
         11550 => x"58",
         11551 => x"7d",
         11552 => x"fd",
         11553 => x"2e",
         11554 => x"b8",
         11555 => x"7a",
         11556 => x"e2",
         11557 => x"e4",
         11558 => x"b8",
         11559 => x"2e",
         11560 => x"78",
         11561 => x"d8",
         11562 => x"c8",
         11563 => x"3d",
         11564 => x"52",
         11565 => x"bd",
         11566 => x"7f",
         11567 => x"5b",
         11568 => x"2e",
         11569 => x"1f",
         11570 => x"81",
         11571 => x"5f",
         11572 => x"f5",
         11573 => x"56",
         11574 => x"81",
         11575 => x"80",
         11576 => x"7e",
         11577 => x"56",
         11578 => x"e6",
         11579 => x"ff",
         11580 => x"59",
         11581 => x"75",
         11582 => x"76",
         11583 => x"18",
         11584 => x"08",
         11585 => x"af",
         11586 => x"da",
         11587 => x"79",
         11588 => x"77",
         11589 => x"8a",
         11590 => x"84",
         11591 => x"70",
         11592 => x"e4",
         11593 => x"08",
         11594 => x"59",
         11595 => x"7e",
         11596 => x"38",
         11597 => x"17",
         11598 => x"5f",
         11599 => x"38",
         11600 => x"7a",
         11601 => x"38",
         11602 => x"7a",
         11603 => x"76",
         11604 => x"33",
         11605 => x"05",
         11606 => x"17",
         11607 => x"26",
         11608 => x"7c",
         11609 => x"5e",
         11610 => x"2e",
         11611 => x"81",
         11612 => x"59",
         11613 => x"78",
         11614 => x"0c",
         11615 => x"0d",
         11616 => x"33",
         11617 => x"71",
         11618 => x"90",
         11619 => x"07",
         11620 => x"fd",
         11621 => x"16",
         11622 => x"33",
         11623 => x"71",
         11624 => x"79",
         11625 => x"3d",
         11626 => x"80",
         11627 => x"ff",
         11628 => x"84",
         11629 => x"59",
         11630 => x"08",
         11631 => x"96",
         11632 => x"39",
         11633 => x"16",
         11634 => x"16",
         11635 => x"17",
         11636 => x"ff",
         11637 => x"81",
         11638 => x"e4",
         11639 => x"38",
         11640 => x"08",
         11641 => x"b4",
         11642 => x"17",
         11643 => x"b8",
         11644 => x"55",
         11645 => x"08",
         11646 => x"38",
         11647 => x"55",
         11648 => x"09",
         11649 => x"f6",
         11650 => x"b4",
         11651 => x"17",
         11652 => x"7d",
         11653 => x"33",
         11654 => x"b8",
         11655 => x"fb",
         11656 => x"18",
         11657 => x"08",
         11658 => x"af",
         11659 => x"0b",
         11660 => x"33",
         11661 => x"83",
         11662 => x"70",
         11663 => x"43",
         11664 => x"5a",
         11665 => x"09",
         11666 => x"e8",
         11667 => x"39",
         11668 => x"08",
         11669 => x"59",
         11670 => x"7c",
         11671 => x"5e",
         11672 => x"27",
         11673 => x"80",
         11674 => x"18",
         11675 => x"5a",
         11676 => x"70",
         11677 => x"34",
         11678 => x"d4",
         11679 => x"39",
         11680 => x"7c",
         11681 => x"b8",
         11682 => x"e4",
         11683 => x"f7",
         11684 => x"7d",
         11685 => x"56",
         11686 => x"9f",
         11687 => x"54",
         11688 => x"97",
         11689 => x"53",
         11690 => x"8f",
         11691 => x"22",
         11692 => x"59",
         11693 => x"2e",
         11694 => x"80",
         11695 => x"75",
         11696 => x"c2",
         11697 => x"33",
         11698 => x"ba",
         11699 => x"08",
         11700 => x"26",
         11701 => x"94",
         11702 => x"80",
         11703 => x"2e",
         11704 => x"79",
         11705 => x"70",
         11706 => x"5a",
         11707 => x"2e",
         11708 => x"75",
         11709 => x"51",
         11710 => x"3f",
         11711 => x"08",
         11712 => x"54",
         11713 => x"53",
         11714 => x"3f",
         11715 => x"08",
         11716 => x"d5",
         11717 => x"74",
         11718 => x"17",
         11719 => x"31",
         11720 => x"56",
         11721 => x"80",
         11722 => x"38",
         11723 => x"81",
         11724 => x"76",
         11725 => x"08",
         11726 => x"0c",
         11727 => x"70",
         11728 => x"06",
         11729 => x"78",
         11730 => x"fe",
         11731 => x"74",
         11732 => x"f3",
         11733 => x"e4",
         11734 => x"b8",
         11735 => x"2e",
         11736 => x"73",
         11737 => x"38",
         11738 => x"82",
         11739 => x"53",
         11740 => x"08",
         11741 => x"38",
         11742 => x"0c",
         11743 => x"81",
         11744 => x"34",
         11745 => x"84",
         11746 => x"8b",
         11747 => x"90",
         11748 => x"81",
         11749 => x"55",
         11750 => x"bb",
         11751 => x"16",
         11752 => x"80",
         11753 => x"2e",
         11754 => x"fe",
         11755 => x"94",
         11756 => x"15",
         11757 => x"74",
         11758 => x"73",
         11759 => x"90",
         11760 => x"c0",
         11761 => x"90",
         11762 => x"83",
         11763 => x"78",
         11764 => x"38",
         11765 => x"78",
         11766 => x"77",
         11767 => x"80",
         11768 => x"e4",
         11769 => x"0d",
         11770 => x"94",
         11771 => x"15",
         11772 => x"80",
         11773 => x"38",
         11774 => x"0c",
         11775 => x"80",
         11776 => x"a8",
         11777 => x"e4",
         11778 => x"15",
         11779 => x"16",
         11780 => x"ff",
         11781 => x"80",
         11782 => x"79",
         11783 => x"12",
         11784 => x"5a",
         11785 => x"78",
         11786 => x"38",
         11787 => x"74",
         11788 => x"18",
         11789 => x"89",
         11790 => x"5a",
         11791 => x"2e",
         11792 => x"8c",
         11793 => x"fe",
         11794 => x"52",
         11795 => x"89",
         11796 => x"b8",
         11797 => x"fe",
         11798 => x"14",
         11799 => x"82",
         11800 => x"b8",
         11801 => x"06",
         11802 => x"cf",
         11803 => x"08",
         11804 => x"c9",
         11805 => x"74",
         11806 => x"cb",
         11807 => x"e4",
         11808 => x"b8",
         11809 => x"2e",
         11810 => x"b8",
         11811 => x"2e",
         11812 => x"84",
         11813 => x"88",
         11814 => x"98",
         11815 => x"dc",
         11816 => x"91",
         11817 => x"0b",
         11818 => x"0c",
         11819 => x"04",
         11820 => x"7c",
         11821 => x"75",
         11822 => x"38",
         11823 => x"3d",
         11824 => x"8d",
         11825 => x"51",
         11826 => x"84",
         11827 => x"55",
         11828 => x"08",
         11829 => x"38",
         11830 => x"74",
         11831 => x"b8",
         11832 => x"3d",
         11833 => x"76",
         11834 => x"75",
         11835 => x"97",
         11836 => x"e4",
         11837 => x"b8",
         11838 => x"d1",
         11839 => x"33",
         11840 => x"59",
         11841 => x"24",
         11842 => x"16",
         11843 => x"2a",
         11844 => x"54",
         11845 => x"80",
         11846 => x"16",
         11847 => x"33",
         11848 => x"71",
         11849 => x"7d",
         11850 => x"5d",
         11851 => x"78",
         11852 => x"38",
         11853 => x"0c",
         11854 => x"18",
         11855 => x"23",
         11856 => x"51",
         11857 => x"3f",
         11858 => x"08",
         11859 => x"2e",
         11860 => x"80",
         11861 => x"38",
         11862 => x"fe",
         11863 => x"55",
         11864 => x"fe",
         11865 => x"17",
         11866 => x"33",
         11867 => x"71",
         11868 => x"7a",
         11869 => x"0c",
         11870 => x"bc",
         11871 => x"0d",
         11872 => x"54",
         11873 => x"9e",
         11874 => x"53",
         11875 => x"96",
         11876 => x"52",
         11877 => x"8e",
         11878 => x"22",
         11879 => x"57",
         11880 => x"2e",
         11881 => x"52",
         11882 => x"84",
         11883 => x"0c",
         11884 => x"e4",
         11885 => x"0d",
         11886 => x"33",
         11887 => x"c3",
         11888 => x"e4",
         11889 => x"52",
         11890 => x"71",
         11891 => x"54",
         11892 => x"3d",
         11893 => x"58",
         11894 => x"74",
         11895 => x"38",
         11896 => x"73",
         11897 => x"38",
         11898 => x"72",
         11899 => x"38",
         11900 => x"84",
         11901 => x"53",
         11902 => x"81",
         11903 => x"53",
         11904 => x"53",
         11905 => x"38",
         11906 => x"80",
         11907 => x"52",
         11908 => x"9d",
         11909 => x"b8",
         11910 => x"84",
         11911 => x"84",
         11912 => x"84",
         11913 => x"a6",
         11914 => x"74",
         11915 => x"92",
         11916 => x"74",
         11917 => x"be",
         11918 => x"e4",
         11919 => x"70",
         11920 => x"07",
         11921 => x"b8",
         11922 => x"55",
         11923 => x"84",
         11924 => x"8a",
         11925 => x"75",
         11926 => x"52",
         11927 => x"e2",
         11928 => x"74",
         11929 => x"8e",
         11930 => x"e4",
         11931 => x"70",
         11932 => x"07",
         11933 => x"b8",
         11934 => x"55",
         11935 => x"39",
         11936 => x"51",
         11937 => x"3f",
         11938 => x"08",
         11939 => x"0c",
         11940 => x"04",
         11941 => x"51",
         11942 => x"3f",
         11943 => x"08",
         11944 => x"72",
         11945 => x"72",
         11946 => x"56",
         11947 => x"ed",
         11948 => x"57",
         11949 => x"3d",
         11950 => x"3d",
         11951 => x"a5",
         11952 => x"e4",
         11953 => x"b8",
         11954 => x"2e",
         11955 => x"84",
         11956 => x"95",
         11957 => x"65",
         11958 => x"ff",
         11959 => x"84",
         11960 => x"55",
         11961 => x"08",
         11962 => x"80",
         11963 => x"70",
         11964 => x"58",
         11965 => x"97",
         11966 => x"2e",
         11967 => x"52",
         11968 => x"b0",
         11969 => x"84",
         11970 => x"95",
         11971 => x"86",
         11972 => x"e4",
         11973 => x"0d",
         11974 => x"0d",
         11975 => x"5f",
         11976 => x"3d",
         11977 => x"96",
         11978 => x"b9",
         11979 => x"e4",
         11980 => x"b8",
         11981 => x"38",
         11982 => x"74",
         11983 => x"08",
         11984 => x"13",
         11985 => x"59",
         11986 => x"26",
         11987 => x"7f",
         11988 => x"b8",
         11989 => x"3d",
         11990 => x"b8",
         11991 => x"33",
         11992 => x"81",
         11993 => x"38",
         11994 => x"08",
         11995 => x"08",
         11996 => x"77",
         11997 => x"7b",
         11998 => x"5c",
         11999 => x"17",
         12000 => x"82",
         12001 => x"17",
         12002 => x"5d",
         12003 => x"38",
         12004 => x"53",
         12005 => x"81",
         12006 => x"fe",
         12007 => x"84",
         12008 => x"80",
         12009 => x"ff",
         12010 => x"79",
         12011 => x"7f",
         12012 => x"7d",
         12013 => x"76",
         12014 => x"82",
         12015 => x"38",
         12016 => x"05",
         12017 => x"82",
         12018 => x"90",
         12019 => x"2b",
         12020 => x"33",
         12021 => x"88",
         12022 => x"71",
         12023 => x"fe",
         12024 => x"70",
         12025 => x"25",
         12026 => x"84",
         12027 => x"06",
         12028 => x"43",
         12029 => x"54",
         12030 => x"40",
         12031 => x"fe",
         12032 => x"7f",
         12033 => x"18",
         12034 => x"33",
         12035 => x"77",
         12036 => x"79",
         12037 => x"0c",
         12038 => x"04",
         12039 => x"17",
         12040 => x"17",
         12041 => x"18",
         12042 => x"fe",
         12043 => x"81",
         12044 => x"e4",
         12045 => x"38",
         12046 => x"08",
         12047 => x"b4",
         12048 => x"18",
         12049 => x"b8",
         12050 => x"55",
         12051 => x"08",
         12052 => x"38",
         12053 => x"55",
         12054 => x"09",
         12055 => x"b0",
         12056 => x"b4",
         12057 => x"18",
         12058 => x"7c",
         12059 => x"33",
         12060 => x"e0",
         12061 => x"fe",
         12062 => x"77",
         12063 => x"59",
         12064 => x"77",
         12065 => x"80",
         12066 => x"e4",
         12067 => x"80",
         12068 => x"b8",
         12069 => x"2e",
         12070 => x"84",
         12071 => x"30",
         12072 => x"e4",
         12073 => x"25",
         12074 => x"18",
         12075 => x"5c",
         12076 => x"08",
         12077 => x"38",
         12078 => x"7a",
         12079 => x"84",
         12080 => x"07",
         12081 => x"18",
         12082 => x"39",
         12083 => x"05",
         12084 => x"71",
         12085 => x"2b",
         12086 => x"70",
         12087 => x"82",
         12088 => x"06",
         12089 => x"5d",
         12090 => x"5f",
         12091 => x"83",
         12092 => x"39",
         12093 => x"bf",
         12094 => x"58",
         12095 => x"0c",
         12096 => x"0c",
         12097 => x"81",
         12098 => x"84",
         12099 => x"83",
         12100 => x"58",
         12101 => x"f7",
         12102 => x"57",
         12103 => x"80",
         12104 => x"76",
         12105 => x"80",
         12106 => x"74",
         12107 => x"80",
         12108 => x"86",
         12109 => x"18",
         12110 => x"78",
         12111 => x"da",
         12112 => x"73",
         12113 => x"dc",
         12114 => x"33",
         12115 => x"d4",
         12116 => x"33",
         12117 => x"81",
         12118 => x"87",
         12119 => x"2e",
         12120 => x"94",
         12121 => x"73",
         12122 => x"27",
         12123 => x"81",
         12124 => x"17",
         12125 => x"57",
         12126 => x"27",
         12127 => x"16",
         12128 => x"b3",
         12129 => x"80",
         12130 => x"0c",
         12131 => x"8c",
         12132 => x"80",
         12133 => x"78",
         12134 => x"75",
         12135 => x"38",
         12136 => x"34",
         12137 => x"84",
         12138 => x"8b",
         12139 => x"78",
         12140 => x"27",
         12141 => x"73",
         12142 => x"fe",
         12143 => x"84",
         12144 => x"59",
         12145 => x"08",
         12146 => x"e9",
         12147 => x"e4",
         12148 => x"82",
         12149 => x"b8",
         12150 => x"2e",
         12151 => x"80",
         12152 => x"75",
         12153 => x"81",
         12154 => x"e4",
         12155 => x"38",
         12156 => x"fe",
         12157 => x"08",
         12158 => x"74",
         12159 => x"af",
         12160 => x"94",
         12161 => x"16",
         12162 => x"54",
         12163 => x"34",
         12164 => x"79",
         12165 => x"38",
         12166 => x"15",
         12167 => x"f6",
         12168 => x"b8",
         12169 => x"06",
         12170 => x"95",
         12171 => x"08",
         12172 => x"8f",
         12173 => x"90",
         12174 => x"54",
         12175 => x"0b",
         12176 => x"fe",
         12177 => x"17",
         12178 => x"51",
         12179 => x"3f",
         12180 => x"08",
         12181 => x"c2",
         12182 => x"e4",
         12183 => x"81",
         12184 => x"81",
         12185 => x"58",
         12186 => x"08",
         12187 => x"27",
         12188 => x"84",
         12189 => x"98",
         12190 => x"08",
         12191 => x"81",
         12192 => x"e4",
         12193 => x"a1",
         12194 => x"e4",
         12195 => x"08",
         12196 => x"38",
         12197 => x"97",
         12198 => x"74",
         12199 => x"ff",
         12200 => x"84",
         12201 => x"55",
         12202 => x"08",
         12203 => x"73",
         12204 => x"fe",
         12205 => x"84",
         12206 => x"59",
         12207 => x"08",
         12208 => x"cb",
         12209 => x"e4",
         12210 => x"80",
         12211 => x"b8",
         12212 => x"2e",
         12213 => x"80",
         12214 => x"75",
         12215 => x"89",
         12216 => x"e4",
         12217 => x"38",
         12218 => x"fe",
         12219 => x"08",
         12220 => x"74",
         12221 => x"38",
         12222 => x"17",
         12223 => x"33",
         12224 => x"73",
         12225 => x"78",
         12226 => x"26",
         12227 => x"80",
         12228 => x"90",
         12229 => x"fc",
         12230 => x"56",
         12231 => x"82",
         12232 => x"33",
         12233 => x"e4",
         12234 => x"e7",
         12235 => x"90",
         12236 => x"54",
         12237 => x"84",
         12238 => x"90",
         12239 => x"54",
         12240 => x"81",
         12241 => x"33",
         12242 => x"f0",
         12243 => x"e4",
         12244 => x"39",
         12245 => x"bb",
         12246 => x"0d",
         12247 => x"3d",
         12248 => x"52",
         12249 => x"ff",
         12250 => x"84",
         12251 => x"56",
         12252 => x"08",
         12253 => x"38",
         12254 => x"e4",
         12255 => x"0d",
         12256 => x"a8",
         12257 => x"9b",
         12258 => x"59",
         12259 => x"3f",
         12260 => x"08",
         12261 => x"e4",
         12262 => x"02",
         12263 => x"33",
         12264 => x"81",
         12265 => x"86",
         12266 => x"38",
         12267 => x"5b",
         12268 => x"c4",
         12269 => x"ee",
         12270 => x"81",
         12271 => x"87",
         12272 => x"b4",
         12273 => x"3d",
         12274 => x"33",
         12275 => x"71",
         12276 => x"73",
         12277 => x"5c",
         12278 => x"83",
         12279 => x"38",
         12280 => x"81",
         12281 => x"80",
         12282 => x"38",
         12283 => x"18",
         12284 => x"ff",
         12285 => x"5f",
         12286 => x"b8",
         12287 => x"8f",
         12288 => x"55",
         12289 => x"3f",
         12290 => x"08",
         12291 => x"e4",
         12292 => x"38",
         12293 => x"08",
         12294 => x"ff",
         12295 => x"84",
         12296 => x"56",
         12297 => x"08",
         12298 => x"0b",
         12299 => x"0c",
         12300 => x"04",
         12301 => x"94",
         12302 => x"98",
         12303 => x"2b",
         12304 => x"5d",
         12305 => x"98",
         12306 => x"e4",
         12307 => x"88",
         12308 => x"e4",
         12309 => x"38",
         12310 => x"a8",
         12311 => x"5d",
         12312 => x"2e",
         12313 => x"74",
         12314 => x"ff",
         12315 => x"84",
         12316 => x"56",
         12317 => x"08",
         12318 => x"38",
         12319 => x"77",
         12320 => x"56",
         12321 => x"2e",
         12322 => x"80",
         12323 => x"7a",
         12324 => x"55",
         12325 => x"89",
         12326 => x"08",
         12327 => x"fd",
         12328 => x"75",
         12329 => x"7d",
         12330 => x"db",
         12331 => x"e4",
         12332 => x"e4",
         12333 => x"0d",
         12334 => x"5d",
         12335 => x"56",
         12336 => x"17",
         12337 => x"82",
         12338 => x"17",
         12339 => x"55",
         12340 => x"09",
         12341 => x"dd",
         12342 => x"75",
         12343 => x"52",
         12344 => x"51",
         12345 => x"3f",
         12346 => x"08",
         12347 => x"38",
         12348 => x"58",
         12349 => x"0c",
         12350 => x"ab",
         12351 => x"08",
         12352 => x"34",
         12353 => x"18",
         12354 => x"08",
         12355 => x"ec",
         12356 => x"78",
         12357 => x"de",
         12358 => x"e4",
         12359 => x"b8",
         12360 => x"2e",
         12361 => x"75",
         12362 => x"81",
         12363 => x"38",
         12364 => x"c8",
         12365 => x"b4",
         12366 => x"7c",
         12367 => x"33",
         12368 => x"90",
         12369 => x"84",
         12370 => x"7a",
         12371 => x"06",
         12372 => x"84",
         12373 => x"83",
         12374 => x"17",
         12375 => x"08",
         12376 => x"e4",
         12377 => x"74",
         12378 => x"27",
         12379 => x"82",
         12380 => x"74",
         12381 => x"81",
         12382 => x"38",
         12383 => x"17",
         12384 => x"08",
         12385 => x"52",
         12386 => x"51",
         12387 => x"3f",
         12388 => x"c5",
         12389 => x"79",
         12390 => x"e1",
         12391 => x"78",
         12392 => x"e4",
         12393 => x"e4",
         12394 => x"b8",
         12395 => x"2e",
         12396 => x"84",
         12397 => x"81",
         12398 => x"38",
         12399 => x"08",
         12400 => x"cb",
         12401 => x"74",
         12402 => x"fe",
         12403 => x"84",
         12404 => x"b3",
         12405 => x"08",
         12406 => x"19",
         12407 => x"58",
         12408 => x"ff",
         12409 => x"16",
         12410 => x"84",
         12411 => x"07",
         12412 => x"18",
         12413 => x"77",
         12414 => x"a1",
         12415 => x"fd",
         12416 => x"56",
         12417 => x"84",
         12418 => x"56",
         12419 => x"81",
         12420 => x"39",
         12421 => x"82",
         12422 => x"ff",
         12423 => x"a0",
         12424 => x"b2",
         12425 => x"b8",
         12426 => x"84",
         12427 => x"80",
         12428 => x"75",
         12429 => x"0c",
         12430 => x"04",
         12431 => x"52",
         12432 => x"52",
         12433 => x"bf",
         12434 => x"e4",
         12435 => x"b8",
         12436 => x"38",
         12437 => x"b8",
         12438 => x"3d",
         12439 => x"b8",
         12440 => x"2e",
         12441 => x"cb",
         12442 => x"f3",
         12443 => x"85",
         12444 => x"56",
         12445 => x"74",
         12446 => x"7d",
         12447 => x"8f",
         12448 => x"5d",
         12449 => x"3f",
         12450 => x"08",
         12451 => x"84",
         12452 => x"83",
         12453 => x"84",
         12454 => x"81",
         12455 => x"38",
         12456 => x"08",
         12457 => x"cb",
         12458 => x"c9",
         12459 => x"b8",
         12460 => x"12",
         12461 => x"57",
         12462 => x"38",
         12463 => x"18",
         12464 => x"5a",
         12465 => x"75",
         12466 => x"38",
         12467 => x"76",
         12468 => x"19",
         12469 => x"58",
         12470 => x"0c",
         12471 => x"84",
         12472 => x"55",
         12473 => x"81",
         12474 => x"ff",
         12475 => x"f4",
         12476 => x"8a",
         12477 => x"77",
         12478 => x"f9",
         12479 => x"77",
         12480 => x"52",
         12481 => x"51",
         12482 => x"3f",
         12483 => x"08",
         12484 => x"81",
         12485 => x"39",
         12486 => x"84",
         12487 => x"b4",
         12488 => x"b8",
         12489 => x"81",
         12490 => x"58",
         12491 => x"3f",
         12492 => x"b8",
         12493 => x"38",
         12494 => x"08",
         12495 => x"b4",
         12496 => x"18",
         12497 => x"74",
         12498 => x"27",
         12499 => x"82",
         12500 => x"7a",
         12501 => x"81",
         12502 => x"38",
         12503 => x"17",
         12504 => x"08",
         12505 => x"52",
         12506 => x"51",
         12507 => x"3f",
         12508 => x"81",
         12509 => x"08",
         12510 => x"7c",
         12511 => x"38",
         12512 => x"08",
         12513 => x"38",
         12514 => x"51",
         12515 => x"3f",
         12516 => x"08",
         12517 => x"e4",
         12518 => x"fd",
         12519 => x"b8",
         12520 => x"2e",
         12521 => x"84",
         12522 => x"ff",
         12523 => x"38",
         12524 => x"52",
         12525 => x"f9",
         12526 => x"b8",
         12527 => x"f3",
         12528 => x"08",
         12529 => x"19",
         12530 => x"59",
         12531 => x"90",
         12532 => x"94",
         12533 => x"17",
         12534 => x"5c",
         12535 => x"34",
         12536 => x"7a",
         12537 => x"38",
         12538 => x"e4",
         12539 => x"0d",
         12540 => x"22",
         12541 => x"ff",
         12542 => x"81",
         12543 => x"2e",
         12544 => x"fe",
         12545 => x"0b",
         12546 => x"56",
         12547 => x"81",
         12548 => x"ff",
         12549 => x"f4",
         12550 => x"ae",
         12551 => x"34",
         12552 => x"0b",
         12553 => x"34",
         12554 => x"80",
         12555 => x"75",
         12556 => x"34",
         12557 => x"d0",
         12558 => x"cc",
         12559 => x"1a",
         12560 => x"83",
         12561 => x"59",
         12562 => x"d2",
         12563 => x"88",
         12564 => x"80",
         12565 => x"75",
         12566 => x"83",
         12567 => x"38",
         12568 => x"0b",
         12569 => x"b8",
         12570 => x"56",
         12571 => x"05",
         12572 => x"70",
         12573 => x"34",
         12574 => x"75",
         12575 => x"56",
         12576 => x"d9",
         12577 => x"7e",
         12578 => x"ff",
         12579 => x"57",
         12580 => x"17",
         12581 => x"2a",
         12582 => x"f3",
         12583 => x"33",
         12584 => x"2e",
         12585 => x"7d",
         12586 => x"83",
         12587 => x"51",
         12588 => x"3f",
         12589 => x"08",
         12590 => x"e4",
         12591 => x"38",
         12592 => x"b8",
         12593 => x"17",
         12594 => x"e4",
         12595 => x"34",
         12596 => x"17",
         12597 => x"0b",
         12598 => x"7d",
         12599 => x"77",
         12600 => x"77",
         12601 => x"78",
         12602 => x"7c",
         12603 => x"83",
         12604 => x"38",
         12605 => x"0b",
         12606 => x"7d",
         12607 => x"83",
         12608 => x"51",
         12609 => x"3f",
         12610 => x"08",
         12611 => x"b8",
         12612 => x"3d",
         12613 => x"90",
         12614 => x"80",
         12615 => x"74",
         12616 => x"76",
         12617 => x"34",
         12618 => x"7b",
         12619 => x"7a",
         12620 => x"34",
         12621 => x"55",
         12622 => x"17",
         12623 => x"a0",
         12624 => x"1a",
         12625 => x"58",
         12626 => x"39",
         12627 => x"58",
         12628 => x"34",
         12629 => x"5c",
         12630 => x"34",
         12631 => x"0b",
         12632 => x"7d",
         12633 => x"83",
         12634 => x"51",
         12635 => x"3f",
         12636 => x"08",
         12637 => x"39",
         12638 => x"b3",
         12639 => x"08",
         12640 => x"5f",
         12641 => x"9b",
         12642 => x"81",
         12643 => x"70",
         12644 => x"56",
         12645 => x"81",
         12646 => x"ed",
         12647 => x"2e",
         12648 => x"82",
         12649 => x"fe",
         12650 => x"b2",
         12651 => x"ab",
         12652 => x"b8",
         12653 => x"84",
         12654 => x"80",
         12655 => x"75",
         12656 => x"0c",
         12657 => x"04",
         12658 => x"0c",
         12659 => x"52",
         12660 => x"52",
         12661 => x"af",
         12662 => x"e4",
         12663 => x"b8",
         12664 => x"38",
         12665 => x"05",
         12666 => x"06",
         12667 => x"7c",
         12668 => x"0b",
         12669 => x"3d",
         12670 => x"55",
         12671 => x"05",
         12672 => x"70",
         12673 => x"34",
         12674 => x"74",
         12675 => x"3d",
         12676 => x"7a",
         12677 => x"75",
         12678 => x"57",
         12679 => x"81",
         12680 => x"ff",
         12681 => x"ef",
         12682 => x"08",
         12683 => x"ff",
         12684 => x"84",
         12685 => x"56",
         12686 => x"08",
         12687 => x"6a",
         12688 => x"2e",
         12689 => x"88",
         12690 => x"e4",
         12691 => x"0d",
         12692 => x"d0",
         12693 => x"ff",
         12694 => x"58",
         12695 => x"91",
         12696 => x"78",
         12697 => x"d0",
         12698 => x"78",
         12699 => x"fa",
         12700 => x"08",
         12701 => x"70",
         12702 => x"5e",
         12703 => x"7a",
         12704 => x"5c",
         12705 => x"81",
         12706 => x"ff",
         12707 => x"58",
         12708 => x"26",
         12709 => x"16",
         12710 => x"06",
         12711 => x"9f",
         12712 => x"99",
         12713 => x"e0",
         12714 => x"ff",
         12715 => x"75",
         12716 => x"2a",
         12717 => x"77",
         12718 => x"06",
         12719 => x"ff",
         12720 => x"7a",
         12721 => x"70",
         12722 => x"2a",
         12723 => x"58",
         12724 => x"2e",
         12725 => x"1c",
         12726 => x"5c",
         12727 => x"fd",
         12728 => x"08",
         12729 => x"ff",
         12730 => x"83",
         12731 => x"38",
         12732 => x"82",
         12733 => x"fe",
         12734 => x"b2",
         12735 => x"a8",
         12736 => x"b8",
         12737 => x"84",
         12738 => x"fd",
         12739 => x"b8",
         12740 => x"3d",
         12741 => x"81",
         12742 => x"38",
         12743 => x"8d",
         12744 => x"b8",
         12745 => x"84",
         12746 => x"fd",
         12747 => x"58",
         12748 => x"19",
         12749 => x"80",
         12750 => x"56",
         12751 => x"81",
         12752 => x"75",
         12753 => x"57",
         12754 => x"5a",
         12755 => x"02",
         12756 => x"33",
         12757 => x"8b",
         12758 => x"84",
         12759 => x"40",
         12760 => x"38",
         12761 => x"57",
         12762 => x"34",
         12763 => x"0b",
         12764 => x"8b",
         12765 => x"84",
         12766 => x"57",
         12767 => x"2e",
         12768 => x"a7",
         12769 => x"2e",
         12770 => x"7f",
         12771 => x"9a",
         12772 => x"88",
         12773 => x"33",
         12774 => x"57",
         12775 => x"82",
         12776 => x"16",
         12777 => x"fe",
         12778 => x"75",
         12779 => x"c7",
         12780 => x"22",
         12781 => x"b0",
         12782 => x"57",
         12783 => x"2e",
         12784 => x"75",
         12785 => x"b4",
         12786 => x"2e",
         12787 => x"17",
         12788 => x"83",
         12789 => x"54",
         12790 => x"17",
         12791 => x"33",
         12792 => x"f1",
         12793 => x"e4",
         12794 => x"85",
         12795 => x"81",
         12796 => x"18",
         12797 => x"7b",
         12798 => x"56",
         12799 => x"bf",
         12800 => x"33",
         12801 => x"2e",
         12802 => x"bb",
         12803 => x"83",
         12804 => x"5d",
         12805 => x"f2",
         12806 => x"88",
         12807 => x"80",
         12808 => x"76",
         12809 => x"83",
         12810 => x"06",
         12811 => x"90",
         12812 => x"80",
         12813 => x"7d",
         12814 => x"75",
         12815 => x"34",
         12816 => x"0b",
         12817 => x"78",
         12818 => x"08",
         12819 => x"57",
         12820 => x"ff",
         12821 => x"74",
         12822 => x"fe",
         12823 => x"84",
         12824 => x"55",
         12825 => x"08",
         12826 => x"b8",
         12827 => x"19",
         12828 => x"5a",
         12829 => x"77",
         12830 => x"83",
         12831 => x"59",
         12832 => x"2e",
         12833 => x"81",
         12834 => x"54",
         12835 => x"16",
         12836 => x"33",
         12837 => x"bd",
         12838 => x"e4",
         12839 => x"85",
         12840 => x"81",
         12841 => x"17",
         12842 => x"77",
         12843 => x"19",
         12844 => x"7a",
         12845 => x"83",
         12846 => x"19",
         12847 => x"a5",
         12848 => x"78",
         12849 => x"ae",
         12850 => x"e4",
         12851 => x"b8",
         12852 => x"2e",
         12853 => x"82",
         12854 => x"2e",
         12855 => x"74",
         12856 => x"db",
         12857 => x"fe",
         12858 => x"84",
         12859 => x"84",
         12860 => x"b1",
         12861 => x"82",
         12862 => x"e4",
         12863 => x"0d",
         12864 => x"33",
         12865 => x"71",
         12866 => x"90",
         12867 => x"07",
         12868 => x"fd",
         12869 => x"b8",
         12870 => x"2e",
         12871 => x"84",
         12872 => x"80",
         12873 => x"38",
         12874 => x"e4",
         12875 => x"0d",
         12876 => x"b4",
         12877 => x"7b",
         12878 => x"33",
         12879 => x"94",
         12880 => x"84",
         12881 => x"7a",
         12882 => x"06",
         12883 => x"84",
         12884 => x"83",
         12885 => x"16",
         12886 => x"08",
         12887 => x"e4",
         12888 => x"74",
         12889 => x"27",
         12890 => x"82",
         12891 => x"7c",
         12892 => x"81",
         12893 => x"38",
         12894 => x"16",
         12895 => x"08",
         12896 => x"52",
         12897 => x"51",
         12898 => x"3f",
         12899 => x"fa",
         12900 => x"b4",
         12901 => x"b8",
         12902 => x"81",
         12903 => x"5b",
         12904 => x"3f",
         12905 => x"b8",
         12906 => x"c9",
         12907 => x"e4",
         12908 => x"34",
         12909 => x"a8",
         12910 => x"84",
         12911 => x"5d",
         12912 => x"18",
         12913 => x"8e",
         12914 => x"33",
         12915 => x"2e",
         12916 => x"fc",
         12917 => x"54",
         12918 => x"a0",
         12919 => x"53",
         12920 => x"17",
         12921 => x"e0",
         12922 => x"5c",
         12923 => x"ec",
         12924 => x"80",
         12925 => x"02",
         12926 => x"e3",
         12927 => x"57",
         12928 => x"3d",
         12929 => x"97",
         12930 => x"a2",
         12931 => x"b8",
         12932 => x"84",
         12933 => x"80",
         12934 => x"75",
         12935 => x"0c",
         12936 => x"04",
         12937 => x"52",
         12938 => x"05",
         12939 => x"d7",
         12940 => x"e4",
         12941 => x"b8",
         12942 => x"38",
         12943 => x"05",
         12944 => x"06",
         12945 => x"73",
         12946 => x"a7",
         12947 => x"09",
         12948 => x"71",
         12949 => x"06",
         12950 => x"57",
         12951 => x"17",
         12952 => x"81",
         12953 => x"34",
         12954 => x"e2",
         12955 => x"b8",
         12956 => x"b8",
         12957 => x"3d",
         12958 => x"3d",
         12959 => x"82",
         12960 => x"cc",
         12961 => x"3d",
         12962 => x"d9",
         12963 => x"e4",
         12964 => x"b8",
         12965 => x"2e",
         12966 => x"84",
         12967 => x"96",
         12968 => x"78",
         12969 => x"96",
         12970 => x"51",
         12971 => x"3f",
         12972 => x"08",
         12973 => x"e4",
         12974 => x"02",
         12975 => x"33",
         12976 => x"56",
         12977 => x"d2",
         12978 => x"18",
         12979 => x"22",
         12980 => x"07",
         12981 => x"76",
         12982 => x"76",
         12983 => x"74",
         12984 => x"76",
         12985 => x"77",
         12986 => x"76",
         12987 => x"73",
         12988 => x"78",
         12989 => x"83",
         12990 => x"51",
         12991 => x"3f",
         12992 => x"08",
         12993 => x"0c",
         12994 => x"04",
         12995 => x"6b",
         12996 => x"80",
         12997 => x"cc",
         12998 => x"3d",
         12999 => x"c5",
         13000 => x"e4",
         13001 => x"e4",
         13002 => x"84",
         13003 => x"07",
         13004 => x"56",
         13005 => x"2e",
         13006 => x"70",
         13007 => x"56",
         13008 => x"38",
         13009 => x"78",
         13010 => x"56",
         13011 => x"2e",
         13012 => x"81",
         13013 => x"5a",
         13014 => x"2e",
         13015 => x"7c",
         13016 => x"58",
         13017 => x"b4",
         13018 => x"2e",
         13019 => x"83",
         13020 => x"5a",
         13021 => x"2e",
         13022 => x"81",
         13023 => x"54",
         13024 => x"16",
         13025 => x"33",
         13026 => x"c9",
         13027 => x"e4",
         13028 => x"85",
         13029 => x"81",
         13030 => x"17",
         13031 => x"78",
         13032 => x"70",
         13033 => x"80",
         13034 => x"83",
         13035 => x"80",
         13036 => x"84",
         13037 => x"a7",
         13038 => x"b8",
         13039 => x"33",
         13040 => x"71",
         13041 => x"88",
         13042 => x"14",
         13043 => x"07",
         13044 => x"33",
         13045 => x"0c",
         13046 => x"57",
         13047 => x"84",
         13048 => x"9a",
         13049 => x"7c",
         13050 => x"80",
         13051 => x"70",
         13052 => x"f4",
         13053 => x"b8",
         13054 => x"84",
         13055 => x"80",
         13056 => x"38",
         13057 => x"09",
         13058 => x"b8",
         13059 => x"34",
         13060 => x"b0",
         13061 => x"b4",
         13062 => x"b8",
         13063 => x"81",
         13064 => x"5b",
         13065 => x"3f",
         13066 => x"b8",
         13067 => x"2e",
         13068 => x"fe",
         13069 => x"b8",
         13070 => x"17",
         13071 => x"08",
         13072 => x"31",
         13073 => x"08",
         13074 => x"a0",
         13075 => x"fe",
         13076 => x"16",
         13077 => x"82",
         13078 => x"06",
         13079 => x"77",
         13080 => x"08",
         13081 => x"05",
         13082 => x"81",
         13083 => x"fe",
         13084 => x"79",
         13085 => x"76",
         13086 => x"52",
         13087 => x"51",
         13088 => x"3f",
         13089 => x"08",
         13090 => x"8d",
         13091 => x"39",
         13092 => x"51",
         13093 => x"3f",
         13094 => x"08",
         13095 => x"e4",
         13096 => x"38",
         13097 => x"08",
         13098 => x"08",
         13099 => x"59",
         13100 => x"19",
         13101 => x"59",
         13102 => x"75",
         13103 => x"59",
         13104 => x"ec",
         13105 => x"1c",
         13106 => x"76",
         13107 => x"2e",
         13108 => x"ff",
         13109 => x"70",
         13110 => x"58",
         13111 => x"ea",
         13112 => x"39",
         13113 => x"ba",
         13114 => x"0d",
         13115 => x"3d",
         13116 => x"52",
         13117 => x"ff",
         13118 => x"84",
         13119 => x"56",
         13120 => x"08",
         13121 => x"8f",
         13122 => x"7d",
         13123 => x"76",
         13124 => x"58",
         13125 => x"55",
         13126 => x"74",
         13127 => x"70",
         13128 => x"ff",
         13129 => x"58",
         13130 => x"27",
         13131 => x"a2",
         13132 => x"5c",
         13133 => x"ff",
         13134 => x"57",
         13135 => x"f5",
         13136 => x"0c",
         13137 => x"ff",
         13138 => x"38",
         13139 => x"95",
         13140 => x"52",
         13141 => x"08",
         13142 => x"3f",
         13143 => x"08",
         13144 => x"06",
         13145 => x"2e",
         13146 => x"83",
         13147 => x"83",
         13148 => x"70",
         13149 => x"5b",
         13150 => x"80",
         13151 => x"38",
         13152 => x"77",
         13153 => x"81",
         13154 => x"70",
         13155 => x"57",
         13156 => x"80",
         13157 => x"74",
         13158 => x"81",
         13159 => x"75",
         13160 => x"59",
         13161 => x"38",
         13162 => x"27",
         13163 => x"79",
         13164 => x"96",
         13165 => x"77",
         13166 => x"76",
         13167 => x"74",
         13168 => x"05",
         13169 => x"1a",
         13170 => x"70",
         13171 => x"34",
         13172 => x"3d",
         13173 => x"70",
         13174 => x"5b",
         13175 => x"77",
         13176 => x"d1",
         13177 => x"33",
         13178 => x"76",
         13179 => x"bc",
         13180 => x"2e",
         13181 => x"b7",
         13182 => x"16",
         13183 => x"5c",
         13184 => x"09",
         13185 => x"38",
         13186 => x"79",
         13187 => x"45",
         13188 => x"52",
         13189 => x"52",
         13190 => x"e4",
         13191 => x"e4",
         13192 => x"b8",
         13193 => x"2e",
         13194 => x"56",
         13195 => x"e4",
         13196 => x"0d",
         13197 => x"52",
         13198 => x"e7",
         13199 => x"e4",
         13200 => x"ff",
         13201 => x"fd",
         13202 => x"56",
         13203 => x"e4",
         13204 => x"0d",
         13205 => x"f4",
         13206 => x"c3",
         13207 => x"75",
         13208 => x"ee",
         13209 => x"e4",
         13210 => x"b8",
         13211 => x"c1",
         13212 => x"2e",
         13213 => x"8b",
         13214 => x"57",
         13215 => x"81",
         13216 => x"76",
         13217 => x"58",
         13218 => x"55",
         13219 => x"7d",
         13220 => x"83",
         13221 => x"51",
         13222 => x"3f",
         13223 => x"08",
         13224 => x"ff",
         13225 => x"7a",
         13226 => x"38",
         13227 => x"9c",
         13228 => x"e4",
         13229 => x"09",
         13230 => x"ee",
         13231 => x"79",
         13232 => x"e6",
         13233 => x"75",
         13234 => x"58",
         13235 => x"3f",
         13236 => x"08",
         13237 => x"e4",
         13238 => x"09",
         13239 => x"84",
         13240 => x"e4",
         13241 => x"5c",
         13242 => x"08",
         13243 => x"b4",
         13244 => x"2e",
         13245 => x"18",
         13246 => x"79",
         13247 => x"06",
         13248 => x"81",
         13249 => x"b8",
         13250 => x"18",
         13251 => x"d5",
         13252 => x"b8",
         13253 => x"2e",
         13254 => x"57",
         13255 => x"b4",
         13256 => x"57",
         13257 => x"78",
         13258 => x"70",
         13259 => x"57",
         13260 => x"2e",
         13261 => x"74",
         13262 => x"25",
         13263 => x"5c",
         13264 => x"81",
         13265 => x"1a",
         13266 => x"2e",
         13267 => x"52",
         13268 => x"ef",
         13269 => x"b8",
         13270 => x"84",
         13271 => x"80",
         13272 => x"38",
         13273 => x"84",
         13274 => x"38",
         13275 => x"fd",
         13276 => x"6c",
         13277 => x"76",
         13278 => x"58",
         13279 => x"55",
         13280 => x"6b",
         13281 => x"8b",
         13282 => x"6c",
         13283 => x"55",
         13284 => x"05",
         13285 => x"70",
         13286 => x"34",
         13287 => x"74",
         13288 => x"eb",
         13289 => x"81",
         13290 => x"76",
         13291 => x"58",
         13292 => x"55",
         13293 => x"fd",
         13294 => x"5a",
         13295 => x"7d",
         13296 => x"83",
         13297 => x"51",
         13298 => x"3f",
         13299 => x"08",
         13300 => x"39",
         13301 => x"df",
         13302 => x"b4",
         13303 => x"7a",
         13304 => x"33",
         13305 => x"ec",
         13306 => x"e4",
         13307 => x"09",
         13308 => x"c3",
         13309 => x"e4",
         13310 => x"34",
         13311 => x"a8",
         13312 => x"5c",
         13313 => x"08",
         13314 => x"82",
         13315 => x"74",
         13316 => x"38",
         13317 => x"08",
         13318 => x"39",
         13319 => x"52",
         13320 => x"ed",
         13321 => x"b8",
         13322 => x"84",
         13323 => x"80",
         13324 => x"38",
         13325 => x"81",
         13326 => x"78",
         13327 => x"e7",
         13328 => x"39",
         13329 => x"18",
         13330 => x"08",
         13331 => x"52",
         13332 => x"51",
         13333 => x"3f",
         13334 => x"f2",
         13335 => x"62",
         13336 => x"80",
         13337 => x"5e",
         13338 => x"56",
         13339 => x"9f",
         13340 => x"55",
         13341 => x"97",
         13342 => x"54",
         13343 => x"8f",
         13344 => x"22",
         13345 => x"59",
         13346 => x"2e",
         13347 => x"80",
         13348 => x"75",
         13349 => x"91",
         13350 => x"75",
         13351 => x"79",
         13352 => x"a2",
         13353 => x"08",
         13354 => x"90",
         13355 => x"81",
         13356 => x"56",
         13357 => x"2e",
         13358 => x"7e",
         13359 => x"70",
         13360 => x"55",
         13361 => x"5c",
         13362 => x"dc",
         13363 => x"7a",
         13364 => x"70",
         13365 => x"2a",
         13366 => x"08",
         13367 => x"08",
         13368 => x"5f",
         13369 => x"78",
         13370 => x"9c",
         13371 => x"26",
         13372 => x"58",
         13373 => x"5b",
         13374 => x"52",
         13375 => x"d8",
         13376 => x"15",
         13377 => x"9c",
         13378 => x"26",
         13379 => x"55",
         13380 => x"08",
         13381 => x"dc",
         13382 => x"e4",
         13383 => x"81",
         13384 => x"b8",
         13385 => x"c5",
         13386 => x"59",
         13387 => x"bb",
         13388 => x"2e",
         13389 => x"c2",
         13390 => x"75",
         13391 => x"b8",
         13392 => x"3d",
         13393 => x"0b",
         13394 => x"0c",
         13395 => x"04",
         13396 => x"51",
         13397 => x"3f",
         13398 => x"08",
         13399 => x"73",
         13400 => x"73",
         13401 => x"56",
         13402 => x"7b",
         13403 => x"8e",
         13404 => x"56",
         13405 => x"2e",
         13406 => x"18",
         13407 => x"2e",
         13408 => x"73",
         13409 => x"7e",
         13410 => x"dd",
         13411 => x"e4",
         13412 => x"b8",
         13413 => x"a3",
         13414 => x"19",
         13415 => x"59",
         13416 => x"38",
         13417 => x"12",
         13418 => x"80",
         13419 => x"38",
         13420 => x"0c",
         13421 => x"0c",
         13422 => x"80",
         13423 => x"7b",
         13424 => x"9c",
         13425 => x"05",
         13426 => x"58",
         13427 => x"26",
         13428 => x"76",
         13429 => x"16",
         13430 => x"33",
         13431 => x"7c",
         13432 => x"75",
         13433 => x"39",
         13434 => x"97",
         13435 => x"80",
         13436 => x"39",
         13437 => x"c5",
         13438 => x"fe",
         13439 => x"1b",
         13440 => x"39",
         13441 => x"08",
         13442 => x"a3",
         13443 => x"3d",
         13444 => x"05",
         13445 => x"33",
         13446 => x"ff",
         13447 => x"08",
         13448 => x"40",
         13449 => x"85",
         13450 => x"70",
         13451 => x"33",
         13452 => x"56",
         13453 => x"2e",
         13454 => x"74",
         13455 => x"ba",
         13456 => x"38",
         13457 => x"33",
         13458 => x"24",
         13459 => x"75",
         13460 => x"d0",
         13461 => x"08",
         13462 => x"80",
         13463 => x"80",
         13464 => x"16",
         13465 => x"11",
         13466 => x"d9",
         13467 => x"5b",
         13468 => x"79",
         13469 => x"a9",
         13470 => x"e4",
         13471 => x"06",
         13472 => x"5d",
         13473 => x"7b",
         13474 => x"75",
         13475 => x"06",
         13476 => x"7f",
         13477 => x"9f",
         13478 => x"53",
         13479 => x"51",
         13480 => x"3f",
         13481 => x"08",
         13482 => x"6d",
         13483 => x"2e",
         13484 => x"74",
         13485 => x"26",
         13486 => x"ff",
         13487 => x"55",
         13488 => x"38",
         13489 => x"88",
         13490 => x"7f",
         13491 => x"38",
         13492 => x"0a",
         13493 => x"38",
         13494 => x"06",
         13495 => x"e7",
         13496 => x"2a",
         13497 => x"89",
         13498 => x"2b",
         13499 => x"47",
         13500 => x"2e",
         13501 => x"65",
         13502 => x"25",
         13503 => x"5f",
         13504 => x"83",
         13505 => x"80",
         13506 => x"38",
         13507 => x"53",
         13508 => x"51",
         13509 => x"3f",
         13510 => x"b8",
         13511 => x"95",
         13512 => x"ff",
         13513 => x"83",
         13514 => x"71",
         13515 => x"59",
         13516 => x"77",
         13517 => x"2e",
         13518 => x"82",
         13519 => x"90",
         13520 => x"83",
         13521 => x"44",
         13522 => x"2e",
         13523 => x"83",
         13524 => x"11",
         13525 => x"33",
         13526 => x"71",
         13527 => x"81",
         13528 => x"72",
         13529 => x"75",
         13530 => x"83",
         13531 => x"11",
         13532 => x"33",
         13533 => x"71",
         13534 => x"81",
         13535 => x"72",
         13536 => x"75",
         13537 => x"5c",
         13538 => x"42",
         13539 => x"a3",
         13540 => x"4e",
         13541 => x"4f",
         13542 => x"78",
         13543 => x"80",
         13544 => x"82",
         13545 => x"57",
         13546 => x"26",
         13547 => x"61",
         13548 => x"81",
         13549 => x"63",
         13550 => x"f9",
         13551 => x"06",
         13552 => x"2e",
         13553 => x"81",
         13554 => x"83",
         13555 => x"6e",
         13556 => x"46",
         13557 => x"62",
         13558 => x"c2",
         13559 => x"38",
         13560 => x"57",
         13561 => x"e6",
         13562 => x"58",
         13563 => x"9d",
         13564 => x"26",
         13565 => x"e6",
         13566 => x"10",
         13567 => x"22",
         13568 => x"74",
         13569 => x"38",
         13570 => x"ee",
         13571 => x"78",
         13572 => x"94",
         13573 => x"e4",
         13574 => x"05",
         13575 => x"e4",
         13576 => x"26",
         13577 => x"0b",
         13578 => x"08",
         13579 => x"e4",
         13580 => x"11",
         13581 => x"05",
         13582 => x"83",
         13583 => x"2a",
         13584 => x"a0",
         13585 => x"7d",
         13586 => x"66",
         13587 => x"70",
         13588 => x"31",
         13589 => x"44",
         13590 => x"89",
         13591 => x"1d",
         13592 => x"29",
         13593 => x"31",
         13594 => x"79",
         13595 => x"38",
         13596 => x"7d",
         13597 => x"70",
         13598 => x"56",
         13599 => x"3f",
         13600 => x"08",
         13601 => x"2e",
         13602 => x"62",
         13603 => x"81",
         13604 => x"38",
         13605 => x"0b",
         13606 => x"08",
         13607 => x"38",
         13608 => x"38",
         13609 => x"74",
         13610 => x"89",
         13611 => x"5b",
         13612 => x"8b",
         13613 => x"b8",
         13614 => x"3d",
         13615 => x"f0",
         13616 => x"4e",
         13617 => x"93",
         13618 => x"e4",
         13619 => x"0d",
         13620 => x"0c",
         13621 => x"d0",
         13622 => x"ff",
         13623 => x"57",
         13624 => x"91",
         13625 => x"77",
         13626 => x"d0",
         13627 => x"77",
         13628 => x"b2",
         13629 => x"83",
         13630 => x"5c",
         13631 => x"57",
         13632 => x"81",
         13633 => x"76",
         13634 => x"58",
         13635 => x"12",
         13636 => x"62",
         13637 => x"38",
         13638 => x"81",
         13639 => x"44",
         13640 => x"45",
         13641 => x"89",
         13642 => x"70",
         13643 => x"59",
         13644 => x"70",
         13645 => x"47",
         13646 => x"09",
         13647 => x"38",
         13648 => x"38",
         13649 => x"70",
         13650 => x"07",
         13651 => x"07",
         13652 => x"7a",
         13653 => x"ce",
         13654 => x"84",
         13655 => x"83",
         13656 => x"98",
         13657 => x"f9",
         13658 => x"3d",
         13659 => x"81",
         13660 => x"fe",
         13661 => x"81",
         13662 => x"e4",
         13663 => x"38",
         13664 => x"77",
         13665 => x"e4",
         13666 => x"75",
         13667 => x"5f",
         13668 => x"57",
         13669 => x"fe",
         13670 => x"7f",
         13671 => x"fb",
         13672 => x"fa",
         13673 => x"83",
         13674 => x"38",
         13675 => x"3d",
         13676 => x"95",
         13677 => x"06",
         13678 => x"67",
         13679 => x"f5",
         13680 => x"70",
         13681 => x"43",
         13682 => x"84",
         13683 => x"9f",
         13684 => x"38",
         13685 => x"77",
         13686 => x"80",
         13687 => x"f5",
         13688 => x"76",
         13689 => x"0c",
         13690 => x"84",
         13691 => x"04",
         13692 => x"81",
         13693 => x"38",
         13694 => x"27",
         13695 => x"81",
         13696 => x"57",
         13697 => x"38",
         13698 => x"57",
         13699 => x"70",
         13700 => x"34",
         13701 => x"74",
         13702 => x"61",
         13703 => x"59",
         13704 => x"70",
         13705 => x"33",
         13706 => x"05",
         13707 => x"15",
         13708 => x"38",
         13709 => x"45",
         13710 => x"82",
         13711 => x"34",
         13712 => x"05",
         13713 => x"ff",
         13714 => x"6a",
         13715 => x"34",
         13716 => x"5c",
         13717 => x"05",
         13718 => x"90",
         13719 => x"83",
         13720 => x"5a",
         13721 => x"91",
         13722 => x"9e",
         13723 => x"49",
         13724 => x"05",
         13725 => x"75",
         13726 => x"26",
         13727 => x"75",
         13728 => x"06",
         13729 => x"93",
         13730 => x"88",
         13731 => x"61",
         13732 => x"f8",
         13733 => x"34",
         13734 => x"05",
         13735 => x"99",
         13736 => x"61",
         13737 => x"80",
         13738 => x"34",
         13739 => x"05",
         13740 => x"2a",
         13741 => x"9d",
         13742 => x"90",
         13743 => x"61",
         13744 => x"7e",
         13745 => x"b8",
         13746 => x"b8",
         13747 => x"9f",
         13748 => x"83",
         13749 => x"38",
         13750 => x"05",
         13751 => x"a8",
         13752 => x"61",
         13753 => x"80",
         13754 => x"05",
         13755 => x"ff",
         13756 => x"74",
         13757 => x"34",
         13758 => x"4b",
         13759 => x"05",
         13760 => x"61",
         13761 => x"a9",
         13762 => x"34",
         13763 => x"05",
         13764 => x"59",
         13765 => x"70",
         13766 => x"33",
         13767 => x"05",
         13768 => x"15",
         13769 => x"38",
         13770 => x"05",
         13771 => x"69",
         13772 => x"ff",
         13773 => x"aa",
         13774 => x"54",
         13775 => x"52",
         13776 => x"c6",
         13777 => x"57",
         13778 => x"08",
         13779 => x"60",
         13780 => x"83",
         13781 => x"38",
         13782 => x"55",
         13783 => x"81",
         13784 => x"ff",
         13785 => x"f4",
         13786 => x"41",
         13787 => x"2e",
         13788 => x"87",
         13789 => x"57",
         13790 => x"83",
         13791 => x"76",
         13792 => x"88",
         13793 => x"55",
         13794 => x"81",
         13795 => x"76",
         13796 => x"78",
         13797 => x"05",
         13798 => x"98",
         13799 => x"64",
         13800 => x"65",
         13801 => x"26",
         13802 => x"59",
         13803 => x"53",
         13804 => x"51",
         13805 => x"3f",
         13806 => x"08",
         13807 => x"84",
         13808 => x"55",
         13809 => x"81",
         13810 => x"ff",
         13811 => x"f4",
         13812 => x"77",
         13813 => x"5b",
         13814 => x"7f",
         13815 => x"7f",
         13816 => x"89",
         13817 => x"62",
         13818 => x"38",
         13819 => x"55",
         13820 => x"83",
         13821 => x"74",
         13822 => x"60",
         13823 => x"fe",
         13824 => x"84",
         13825 => x"85",
         13826 => x"1b",
         13827 => x"57",
         13828 => x"38",
         13829 => x"83",
         13830 => x"86",
         13831 => x"ff",
         13832 => x"38",
         13833 => x"82",
         13834 => x"81",
         13835 => x"c1",
         13836 => x"2a",
         13837 => x"7d",
         13838 => x"84",
         13839 => x"59",
         13840 => x"81",
         13841 => x"ff",
         13842 => x"f4",
         13843 => x"69",
         13844 => x"6b",
         13845 => x"be",
         13846 => x"67",
         13847 => x"81",
         13848 => x"67",
         13849 => x"78",
         13850 => x"34",
         13851 => x"05",
         13852 => x"80",
         13853 => x"62",
         13854 => x"f8",
         13855 => x"67",
         13856 => x"84",
         13857 => x"82",
         13858 => x"57",
         13859 => x"05",
         13860 => x"e4",
         13861 => x"05",
         13862 => x"83",
         13863 => x"67",
         13864 => x"05",
         13865 => x"83",
         13866 => x"84",
         13867 => x"61",
         13868 => x"34",
         13869 => x"ca",
         13870 => x"88",
         13871 => x"61",
         13872 => x"34",
         13873 => x"58",
         13874 => x"cc",
         13875 => x"98",
         13876 => x"61",
         13877 => x"34",
         13878 => x"53",
         13879 => x"51",
         13880 => x"3f",
         13881 => x"b8",
         13882 => x"c9",
         13883 => x"80",
         13884 => x"fe",
         13885 => x"81",
         13886 => x"e4",
         13887 => x"38",
         13888 => x"08",
         13889 => x"0c",
         13890 => x"84",
         13891 => x"04",
         13892 => x"e4",
         13893 => x"64",
         13894 => x"f6",
         13895 => x"ae",
         13896 => x"2a",
         13897 => x"83",
         13898 => x"56",
         13899 => x"2e",
         13900 => x"77",
         13901 => x"83",
         13902 => x"77",
         13903 => x"70",
         13904 => x"58",
         13905 => x"86",
         13906 => x"27",
         13907 => x"52",
         13908 => x"f6",
         13909 => x"b8",
         13910 => x"10",
         13911 => x"70",
         13912 => x"5c",
         13913 => x"0b",
         13914 => x"08",
         13915 => x"05",
         13916 => x"ff",
         13917 => x"27",
         13918 => x"8e",
         13919 => x"39",
         13920 => x"08",
         13921 => x"26",
         13922 => x"7a",
         13923 => x"77",
         13924 => x"7a",
         13925 => x"8e",
         13926 => x"39",
         13927 => x"44",
         13928 => x"f8",
         13929 => x"43",
         13930 => x"75",
         13931 => x"34",
         13932 => x"49",
         13933 => x"05",
         13934 => x"2a",
         13935 => x"a2",
         13936 => x"98",
         13937 => x"61",
         13938 => x"f9",
         13939 => x"61",
         13940 => x"34",
         13941 => x"c4",
         13942 => x"61",
         13943 => x"34",
         13944 => x"80",
         13945 => x"7c",
         13946 => x"34",
         13947 => x"5c",
         13948 => x"05",
         13949 => x"2a",
         13950 => x"a6",
         13951 => x"98",
         13952 => x"61",
         13953 => x"82",
         13954 => x"34",
         13955 => x"05",
         13956 => x"ae",
         13957 => x"61",
         13958 => x"81",
         13959 => x"34",
         13960 => x"05",
         13961 => x"b2",
         13962 => x"61",
         13963 => x"ff",
         13964 => x"c0",
         13965 => x"61",
         13966 => x"34",
         13967 => x"c7",
         13968 => x"c0",
         13969 => x"76",
         13970 => x"58",
         13971 => x"81",
         13972 => x"ff",
         13973 => x"80",
         13974 => x"38",
         13975 => x"05",
         13976 => x"70",
         13977 => x"34",
         13978 => x"74",
         13979 => x"b8",
         13980 => x"80",
         13981 => x"79",
         13982 => x"d9",
         13983 => x"84",
         13984 => x"f4",
         13985 => x"90",
         13986 => x"42",
         13987 => x"b2",
         13988 => x"54",
         13989 => x"08",
         13990 => x"79",
         13991 => x"b4",
         13992 => x"39",
         13993 => x"b8",
         13994 => x"3d",
         13995 => x"f0",
         13996 => x"61",
         13997 => x"ff",
         13998 => x"05",
         13999 => x"6a",
         14000 => x"4c",
         14001 => x"34",
         14002 => x"05",
         14003 => x"85",
         14004 => x"61",
         14005 => x"ff",
         14006 => x"34",
         14007 => x"05",
         14008 => x"89",
         14009 => x"61",
         14010 => x"8f",
         14011 => x"57",
         14012 => x"76",
         14013 => x"53",
         14014 => x"51",
         14015 => x"3f",
         14016 => x"56",
         14017 => x"70",
         14018 => x"34",
         14019 => x"76",
         14020 => x"5c",
         14021 => x"70",
         14022 => x"34",
         14023 => x"d2",
         14024 => x"05",
         14025 => x"e1",
         14026 => x"05",
         14027 => x"c1",
         14028 => x"f2",
         14029 => x"05",
         14030 => x"61",
         14031 => x"34",
         14032 => x"83",
         14033 => x"80",
         14034 => x"e7",
         14035 => x"ff",
         14036 => x"61",
         14037 => x"34",
         14038 => x"59",
         14039 => x"e9",
         14040 => x"90",
         14041 => x"61",
         14042 => x"34",
         14043 => x"40",
         14044 => x"eb",
         14045 => x"61",
         14046 => x"34",
         14047 => x"ed",
         14048 => x"61",
         14049 => x"34",
         14050 => x"ef",
         14051 => x"d5",
         14052 => x"aa",
         14053 => x"54",
         14054 => x"60",
         14055 => x"fe",
         14056 => x"81",
         14057 => x"53",
         14058 => x"51",
         14059 => x"3f",
         14060 => x"55",
         14061 => x"f4",
         14062 => x"61",
         14063 => x"7b",
         14064 => x"5a",
         14065 => x"78",
         14066 => x"8d",
         14067 => x"3d",
         14068 => x"81",
         14069 => x"79",
         14070 => x"b4",
         14071 => x"2e",
         14072 => x"9e",
         14073 => x"33",
         14074 => x"2e",
         14075 => x"76",
         14076 => x"58",
         14077 => x"57",
         14078 => x"86",
         14079 => x"24",
         14080 => x"76",
         14081 => x"76",
         14082 => x"55",
         14083 => x"e4",
         14084 => x"0d",
         14085 => x"0d",
         14086 => x"05",
         14087 => x"59",
         14088 => x"2e",
         14089 => x"84",
         14090 => x"80",
         14091 => x"38",
         14092 => x"77",
         14093 => x"56",
         14094 => x"34",
         14095 => x"74",
         14096 => x"38",
         14097 => x"0c",
         14098 => x"18",
         14099 => x"0d",
         14100 => x"fc",
         14101 => x"53",
         14102 => x"76",
         14103 => x"9e",
         14104 => x"7a",
         14105 => x"70",
         14106 => x"2a",
         14107 => x"1b",
         14108 => x"88",
         14109 => x"56",
         14110 => x"8d",
         14111 => x"ff",
         14112 => x"a3",
         14113 => x"0d",
         14114 => x"05",
         14115 => x"58",
         14116 => x"77",
         14117 => x"76",
         14118 => x"58",
         14119 => x"55",
         14120 => x"a1",
         14121 => x"0c",
         14122 => x"80",
         14123 => x"56",
         14124 => x"80",
         14125 => x"77",
         14126 => x"56",
         14127 => x"34",
         14128 => x"74",
         14129 => x"38",
         14130 => x"0c",
         14131 => x"18",
         14132 => x"80",
         14133 => x"38",
         14134 => x"ac",
         14135 => x"54",
         14136 => x"76",
         14137 => x"9d",
         14138 => x"b8",
         14139 => x"38",
         14140 => x"ba",
         14141 => x"84",
         14142 => x"9f",
         14143 => x"9f",
         14144 => x"11",
         14145 => x"c0",
         14146 => x"08",
         14147 => x"a2",
         14148 => x"32",
         14149 => x"72",
         14150 => x"70",
         14151 => x"56",
         14152 => x"39",
         14153 => x"51",
         14154 => x"ff",
         14155 => x"84",
         14156 => x"9f",
         14157 => x"fd",
         14158 => x"02",
         14159 => x"05",
         14160 => x"80",
         14161 => x"ff",
         14162 => x"72",
         14163 => x"06",
         14164 => x"b8",
         14165 => x"3d",
         14166 => x"ff",
         14167 => x"54",
         14168 => x"2e",
         14169 => x"e9",
         14170 => x"2e",
         14171 => x"e6",
         14172 => x"72",
         14173 => x"38",
         14174 => x"83",
         14175 => x"53",
         14176 => x"ff",
         14177 => x"71",
         14178 => x"a8",
         14179 => x"51",
         14180 => x"81",
         14181 => x"81",
         14182 => x"b8",
         14183 => x"85",
         14184 => x"fe",
         14185 => x"92",
         14186 => x"84",
         14187 => x"22",
         14188 => x"53",
         14189 => x"26",
         14190 => x"53",
         14191 => x"e4",
         14192 => x"0d",
         14193 => x"b5",
         14194 => x"06",
         14195 => x"81",
         14196 => x"38",
         14197 => x"e4",
         14198 => x"22",
         14199 => x"0c",
         14200 => x"0d",
         14201 => x"0d",
         14202 => x"83",
         14203 => x"80",
         14204 => x"83",
         14205 => x"83",
         14206 => x"56",
         14207 => x"26",
         14208 => x"74",
         14209 => x"56",
         14210 => x"30",
         14211 => x"73",
         14212 => x"54",
         14213 => x"70",
         14214 => x"70",
         14215 => x"22",
         14216 => x"2a",
         14217 => x"ff",
         14218 => x"52",
         14219 => x"24",
         14220 => x"cf",
         14221 => x"15",
         14222 => x"05",
         14223 => x"73",
         14224 => x"25",
         14225 => x"07",
         14226 => x"70",
         14227 => x"38",
         14228 => x"84",
         14229 => x"87",
         14230 => x"83",
         14231 => x"ff",
         14232 => x"88",
         14233 => x"71",
         14234 => x"c9",
         14235 => x"73",
         14236 => x"a0",
         14237 => x"ff",
         14238 => x"51",
         14239 => x"39",
         14240 => x"70",
         14241 => x"06",
         14242 => x"39",
         14243 => x"83",
         14244 => x"57",
         14245 => x"e6",
         14246 => x"ff",
         14247 => x"51",
         14248 => x"16",
         14249 => x"ff",
         14250 => x"d0",
         14251 => x"70",
         14252 => x"06",
         14253 => x"39",
         14254 => x"83",
         14255 => x"57",
         14256 => x"39",
         14257 => x"81",
         14258 => x"31",
         14259 => x"ff",
         14260 => x"55",
         14261 => x"75",
         14262 => x"75",
         14263 => x"52",
         14264 => x"39",
         14265 => x"00",
         14266 => x"ff",
         14267 => x"ff",
         14268 => x"ff",
         14269 => x"00",
         14270 => x"00",
         14271 => x"00",
         14272 => x"00",
         14273 => x"00",
         14274 => x"00",
         14275 => x"00",
         14276 => x"00",
         14277 => x"00",
         14278 => x"00",
         14279 => x"00",
         14280 => x"00",
         14281 => x"00",
         14282 => x"00",
         14283 => x"00",
         14284 => x"00",
         14285 => x"00",
         14286 => x"00",
         14287 => x"00",
         14288 => x"00",
         14289 => x"00",
         14290 => x"00",
         14291 => x"00",
         14292 => x"00",
         14293 => x"00",
         14294 => x"00",
         14295 => x"00",
         14296 => x"00",
         14297 => x"00",
         14298 => x"00",
         14299 => x"00",
         14300 => x"00",
         14301 => x"00",
         14302 => x"00",
         14303 => x"00",
         14304 => x"00",
         14305 => x"00",
         14306 => x"00",
         14307 => x"00",
         14308 => x"00",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"64",
         14743 => x"74",
         14744 => x"64",
         14745 => x"74",
         14746 => x"66",
         14747 => x"74",
         14748 => x"66",
         14749 => x"64",
         14750 => x"66",
         14751 => x"63",
         14752 => x"6d",
         14753 => x"61",
         14754 => x"6d",
         14755 => x"79",
         14756 => x"6d",
         14757 => x"66",
         14758 => x"6d",
         14759 => x"70",
         14760 => x"6d",
         14761 => x"6d",
         14762 => x"6d",
         14763 => x"68",
         14764 => x"68",
         14765 => x"68",
         14766 => x"68",
         14767 => x"63",
         14768 => x"00",
         14769 => x"6a",
         14770 => x"72",
         14771 => x"61",
         14772 => x"72",
         14773 => x"74",
         14774 => x"69",
         14775 => x"00",
         14776 => x"74",
         14777 => x"00",
         14778 => x"63",
         14779 => x"7a",
         14780 => x"74",
         14781 => x"69",
         14782 => x"6d",
         14783 => x"69",
         14784 => x"6b",
         14785 => x"00",
         14786 => x"65",
         14787 => x"55",
         14788 => x"6f",
         14789 => x"65",
         14790 => x"72",
         14791 => x"50",
         14792 => x"6d",
         14793 => x"72",
         14794 => x"6e",
         14795 => x"72",
         14796 => x"2e",
         14797 => x"54",
         14798 => x"6d",
         14799 => x"20",
         14800 => x"6e",
         14801 => x"6c",
         14802 => x"00",
         14803 => x"49",
         14804 => x"66",
         14805 => x"69",
         14806 => x"20",
         14807 => x"6f",
         14808 => x"00",
         14809 => x"46",
         14810 => x"20",
         14811 => x"6c",
         14812 => x"65",
         14813 => x"54",
         14814 => x"6f",
         14815 => x"20",
         14816 => x"72",
         14817 => x"6f",
         14818 => x"61",
         14819 => x"6c",
         14820 => x"2e",
         14821 => x"46",
         14822 => x"61",
         14823 => x"62",
         14824 => x"65",
         14825 => x"4e",
         14826 => x"6f",
         14827 => x"74",
         14828 => x"65",
         14829 => x"6c",
         14830 => x"73",
         14831 => x"20",
         14832 => x"6e",
         14833 => x"6e",
         14834 => x"73",
         14835 => x"44",
         14836 => x"20",
         14837 => x"20",
         14838 => x"62",
         14839 => x"2e",
         14840 => x"44",
         14841 => x"65",
         14842 => x"6d",
         14843 => x"20",
         14844 => x"69",
         14845 => x"6c",
         14846 => x"00",
         14847 => x"53",
         14848 => x"73",
         14849 => x"69",
         14850 => x"70",
         14851 => x"65",
         14852 => x"64",
         14853 => x"46",
         14854 => x"20",
         14855 => x"64",
         14856 => x"69",
         14857 => x"6c",
         14858 => x"00",
         14859 => x"46",
         14860 => x"20",
         14861 => x"65",
         14862 => x"20",
         14863 => x"73",
         14864 => x"00",
         14865 => x"41",
         14866 => x"73",
         14867 => x"65",
         14868 => x"64",
         14869 => x"49",
         14870 => x"6c",
         14871 => x"66",
         14872 => x"6e",
         14873 => x"2e",
         14874 => x"4e",
         14875 => x"61",
         14876 => x"66",
         14877 => x"64",
         14878 => x"4e",
         14879 => x"69",
         14880 => x"66",
         14881 => x"64",
         14882 => x"44",
         14883 => x"20",
         14884 => x"20",
         14885 => x"64",
         14886 => x"49",
         14887 => x"72",
         14888 => x"20",
         14889 => x"6f",
         14890 => x"44",
         14891 => x"20",
         14892 => x"6f",
         14893 => x"53",
         14894 => x"65",
         14895 => x"00",
         14896 => x"0a",
         14897 => x"20",
         14898 => x"65",
         14899 => x"73",
         14900 => x"20",
         14901 => x"20",
         14902 => x"65",
         14903 => x"65",
         14904 => x"00",
         14905 => x"72",
         14906 => x"00",
         14907 => x"25",
         14908 => x"58",
         14909 => x"3a",
         14910 => x"25",
         14911 => x"00",
         14912 => x"20",
         14913 => x"7c",
         14914 => x"20",
         14915 => x"25",
         14916 => x"00",
         14917 => x"20",
         14918 => x"20",
         14919 => x"00",
         14920 => x"7a",
         14921 => x"2a",
         14922 => x"73",
         14923 => x"31",
         14924 => x"34",
         14925 => x"32",
         14926 => x"76",
         14927 => x"00",
         14928 => x"20",
         14929 => x"2c",
         14930 => x"76",
         14931 => x"32",
         14932 => x"25",
         14933 => x"73",
         14934 => x"0a",
         14935 => x"5a",
         14936 => x"49",
         14937 => x"72",
         14938 => x"74",
         14939 => x"6e",
         14940 => x"72",
         14941 => x"55",
         14942 => x"31",
         14943 => x"20",
         14944 => x"65",
         14945 => x"70",
         14946 => x"55",
         14947 => x"31",
         14948 => x"20",
         14949 => x"65",
         14950 => x"70",
         14951 => x"55",
         14952 => x"30",
         14953 => x"20",
         14954 => x"65",
         14955 => x"70",
         14956 => x"55",
         14957 => x"30",
         14958 => x"20",
         14959 => x"65",
         14960 => x"70",
         14961 => x"49",
         14962 => x"4c",
         14963 => x"20",
         14964 => x"65",
         14965 => x"70",
         14966 => x"49",
         14967 => x"4c",
         14968 => x"20",
         14969 => x"65",
         14970 => x"70",
         14971 => x"50",
         14972 => x"69",
         14973 => x"72",
         14974 => x"74",
         14975 => x"54",
         14976 => x"72",
         14977 => x"74",
         14978 => x"75",
         14979 => x"53",
         14980 => x"69",
         14981 => x"75",
         14982 => x"69",
         14983 => x"2e",
         14984 => x"45",
         14985 => x"6c",
         14986 => x"20",
         14987 => x"65",
         14988 => x"2e",
         14989 => x"61",
         14990 => x"65",
         14991 => x"2e",
         14992 => x"00",
         14993 => x"7a",
         14994 => x"7a",
         14995 => x"68",
         14996 => x"46",
         14997 => x"65",
         14998 => x"6f",
         14999 => x"69",
         15000 => x"6c",
         15001 => x"20",
         15002 => x"63",
         15003 => x"20",
         15004 => x"70",
         15005 => x"73",
         15006 => x"6e",
         15007 => x"6d",
         15008 => x"61",
         15009 => x"2e",
         15010 => x"2a",
         15011 => x"25",
         15012 => x"25",
         15013 => x"30",
         15014 => x"42",
         15015 => x"63",
         15016 => x"61",
         15017 => x"00",
         15018 => x"5a",
         15019 => x"62",
         15020 => x"25",
         15021 => x"25",
         15022 => x"73",
         15023 => x"00",
         15024 => x"43",
         15025 => x"20",
         15026 => x"6f",
         15027 => x"6e",
         15028 => x"2e",
         15029 => x"52",
         15030 => x"61",
         15031 => x"6e",
         15032 => x"70",
         15033 => x"63",
         15034 => x"6f",
         15035 => x"2e",
         15036 => x"43",
         15037 => x"69",
         15038 => x"63",
         15039 => x"20",
         15040 => x"30",
         15041 => x"20",
         15042 => x"0a",
         15043 => x"43",
         15044 => x"20",
         15045 => x"75",
         15046 => x"64",
         15047 => x"64",
         15048 => x"25",
         15049 => x"0a",
         15050 => x"45",
         15051 => x"75",
         15052 => x"67",
         15053 => x"64",
         15054 => x"20",
         15055 => x"6c",
         15056 => x"2e",
         15057 => x"25",
         15058 => x"58",
         15059 => x"38",
         15060 => x"00",
         15061 => x"25",
         15062 => x"58",
         15063 => x"34",
         15064 => x"43",
         15065 => x"61",
         15066 => x"67",
         15067 => x"00",
         15068 => x"25",
         15069 => x"78",
         15070 => x"38",
         15071 => x"3e",
         15072 => x"6c",
         15073 => x"30",
         15074 => x"0a",
         15075 => x"43",
         15076 => x"69",
         15077 => x"2e",
         15078 => x"25",
         15079 => x"58",
         15080 => x"32",
         15081 => x"43",
         15082 => x"72",
         15083 => x"2e",
         15084 => x"00",
         15085 => x"44",
         15086 => x"20",
         15087 => x"6f",
         15088 => x"0a",
         15089 => x"70",
         15090 => x"65",
         15091 => x"25",
         15092 => x"25",
         15093 => x"73",
         15094 => x"4d",
         15095 => x"72",
         15096 => x"78",
         15097 => x"73",
         15098 => x"2c",
         15099 => x"6e",
         15100 => x"20",
         15101 => x"63",
         15102 => x"20",
         15103 => x"6d",
         15104 => x"2e",
         15105 => x"3f",
         15106 => x"25",
         15107 => x"64",
         15108 => x"20",
         15109 => x"25",
         15110 => x"64",
         15111 => x"25",
         15112 => x"53",
         15113 => x"43",
         15114 => x"69",
         15115 => x"61",
         15116 => x"6e",
         15117 => x"3a",
         15118 => x"76",
         15119 => x"73",
         15120 => x"70",
         15121 => x"65",
         15122 => x"64",
         15123 => x"41",
         15124 => x"65",
         15125 => x"73",
         15126 => x"20",
         15127 => x"43",
         15128 => x"52",
         15129 => x"74",
         15130 => x"63",
         15131 => x"20",
         15132 => x"72",
         15133 => x"20",
         15134 => x"30",
         15135 => x"00",
         15136 => x"20",
         15137 => x"43",
         15138 => x"4d",
         15139 => x"72",
         15140 => x"74",
         15141 => x"20",
         15142 => x"72",
         15143 => x"20",
         15144 => x"30",
         15145 => x"00",
         15146 => x"20",
         15147 => x"53",
         15148 => x"6b",
         15149 => x"61",
         15150 => x"41",
         15151 => x"65",
         15152 => x"20",
         15153 => x"20",
         15154 => x"30",
         15155 => x"00",
         15156 => x"4d",
         15157 => x"3a",
         15158 => x"20",
         15159 => x"5a",
         15160 => x"49",
         15161 => x"20",
         15162 => x"20",
         15163 => x"20",
         15164 => x"20",
         15165 => x"20",
         15166 => x"30",
         15167 => x"00",
         15168 => x"20",
         15169 => x"53",
         15170 => x"65",
         15171 => x"6c",
         15172 => x"20",
         15173 => x"71",
         15174 => x"20",
         15175 => x"20",
         15176 => x"64",
         15177 => x"34",
         15178 => x"7a",
         15179 => x"20",
         15180 => x"57",
         15181 => x"62",
         15182 => x"20",
         15183 => x"41",
         15184 => x"6c",
         15185 => x"20",
         15186 => x"71",
         15187 => x"64",
         15188 => x"34",
         15189 => x"7a",
         15190 => x"20",
         15191 => x"53",
         15192 => x"4d",
         15193 => x"6f",
         15194 => x"46",
         15195 => x"20",
         15196 => x"20",
         15197 => x"20",
         15198 => x"64",
         15199 => x"34",
         15200 => x"7a",
         15201 => x"20",
         15202 => x"53",
         15203 => x"20",
         15204 => x"50",
         15205 => x"20",
         15206 => x"49",
         15207 => x"4c",
         15208 => x"20",
         15209 => x"57",
         15210 => x"32",
         15211 => x"20",
         15212 => x"57",
         15213 => x"42",
         15214 => x"20",
         15215 => x"00",
         15216 => x"20",
         15217 => x"49",
         15218 => x"20",
         15219 => x"4c",
         15220 => x"68",
         15221 => x"65",
         15222 => x"25",
         15223 => x"29",
         15224 => x"20",
         15225 => x"54",
         15226 => x"52",
         15227 => x"20",
         15228 => x"69",
         15229 => x"73",
         15230 => x"25",
         15231 => x"29",
         15232 => x"20",
         15233 => x"53",
         15234 => x"41",
         15235 => x"20",
         15236 => x"65",
         15237 => x"65",
         15238 => x"25",
         15239 => x"29",
         15240 => x"20",
         15241 => x"52",
         15242 => x"20",
         15243 => x"20",
         15244 => x"30",
         15245 => x"25",
         15246 => x"29",
         15247 => x"20",
         15248 => x"42",
         15249 => x"20",
         15250 => x"20",
         15251 => x"30",
         15252 => x"25",
         15253 => x"29",
         15254 => x"20",
         15255 => x"49",
         15256 => x"20",
         15257 => x"4d",
         15258 => x"30",
         15259 => x"25",
         15260 => x"29",
         15261 => x"20",
         15262 => x"53",
         15263 => x"4d",
         15264 => x"20",
         15265 => x"30",
         15266 => x"25",
         15267 => x"29",
         15268 => x"20",
         15269 => x"57",
         15270 => x"44",
         15271 => x"20",
         15272 => x"30",
         15273 => x"25",
         15274 => x"29",
         15275 => x"20",
         15276 => x"6f",
         15277 => x"6f",
         15278 => x"6f",
         15279 => x"67",
         15280 => x"55",
         15281 => x"6f",
         15282 => x"45",
         15283 => x"00",
         15284 => x"53",
         15285 => x"6c",
         15286 => x"4d",
         15287 => x"75",
         15288 => x"46",
         15289 => x"00",
         15290 => x"45",
         15291 => x"00",
         15292 => x"01",
         15293 => x"00",
         15294 => x"00",
         15295 => x"01",
         15296 => x"00",
         15297 => x"00",
         15298 => x"01",
         15299 => x"00",
         15300 => x"00",
         15301 => x"01",
         15302 => x"00",
         15303 => x"00",
         15304 => x"01",
         15305 => x"00",
         15306 => x"00",
         15307 => x"01",
         15308 => x"00",
         15309 => x"00",
         15310 => x"01",
         15311 => x"00",
         15312 => x"00",
         15313 => x"01",
         15314 => x"00",
         15315 => x"00",
         15316 => x"01",
         15317 => x"00",
         15318 => x"00",
         15319 => x"01",
         15320 => x"00",
         15321 => x"00",
         15322 => x"01",
         15323 => x"00",
         15324 => x"00",
         15325 => x"04",
         15326 => x"00",
         15327 => x"00",
         15328 => x"04",
         15329 => x"00",
         15330 => x"00",
         15331 => x"04",
         15332 => x"00",
         15333 => x"00",
         15334 => x"03",
         15335 => x"00",
         15336 => x"00",
         15337 => x"04",
         15338 => x"00",
         15339 => x"00",
         15340 => x"04",
         15341 => x"00",
         15342 => x"00",
         15343 => x"04",
         15344 => x"00",
         15345 => x"00",
         15346 => x"03",
         15347 => x"00",
         15348 => x"00",
         15349 => x"03",
         15350 => x"00",
         15351 => x"00",
         15352 => x"03",
         15353 => x"00",
         15354 => x"00",
         15355 => x"03",
         15356 => x"00",
         15357 => x"1b",
         15358 => x"1b",
         15359 => x"1b",
         15360 => x"1b",
         15361 => x"1b",
         15362 => x"1b",
         15363 => x"1b",
         15364 => x"1b",
         15365 => x"1b",
         15366 => x"1b",
         15367 => x"1b",
         15368 => x"10",
         15369 => x"0e",
         15370 => x"0d",
         15371 => x"0b",
         15372 => x"08",
         15373 => x"06",
         15374 => x"05",
         15375 => x"04",
         15376 => x"03",
         15377 => x"02",
         15378 => x"01",
         15379 => x"43",
         15380 => x"6f",
         15381 => x"70",
         15382 => x"63",
         15383 => x"74",
         15384 => x"69",
         15385 => x"72",
         15386 => x"69",
         15387 => x"20",
         15388 => x"61",
         15389 => x"6e",
         15390 => x"68",
         15391 => x"6f",
         15392 => x"68",
         15393 => x"00",
         15394 => x"21",
         15395 => x"25",
         15396 => x"75",
         15397 => x"73",
         15398 => x"46",
         15399 => x"65",
         15400 => x"6f",
         15401 => x"73",
         15402 => x"74",
         15403 => x"68",
         15404 => x"6f",
         15405 => x"66",
         15406 => x"20",
         15407 => x"45",
         15408 => x"00",
         15409 => x"3e",
         15410 => x"00",
         15411 => x"1b",
         15412 => x"00",
         15413 => x"1b",
         15414 => x"1b",
         15415 => x"1b",
         15416 => x"1b",
         15417 => x"1b",
         15418 => x"7e",
         15419 => x"1b",
         15420 => x"7e",
         15421 => x"1b",
         15422 => x"7e",
         15423 => x"1b",
         15424 => x"7e",
         15425 => x"1b",
         15426 => x"7e",
         15427 => x"1b",
         15428 => x"7e",
         15429 => x"1b",
         15430 => x"7e",
         15431 => x"1b",
         15432 => x"7e",
         15433 => x"1b",
         15434 => x"7e",
         15435 => x"1b",
         15436 => x"7e",
         15437 => x"1b",
         15438 => x"00",
         15439 => x"1b",
         15440 => x"00",
         15441 => x"1b",
         15442 => x"1b",
         15443 => x"00",
         15444 => x"1b",
         15445 => x"00",
         15446 => x"58",
         15447 => x"2c",
         15448 => x"25",
         15449 => x"64",
         15450 => x"2c",
         15451 => x"25",
         15452 => x"00",
         15453 => x"44",
         15454 => x"2d",
         15455 => x"25",
         15456 => x"63",
         15457 => x"2c",
         15458 => x"25",
         15459 => x"25",
         15460 => x"4b",
         15461 => x"3a",
         15462 => x"25",
         15463 => x"2c",
         15464 => x"25",
         15465 => x"64",
         15466 => x"52",
         15467 => x"52",
         15468 => x"72",
         15469 => x"75",
         15470 => x"72",
         15471 => x"55",
         15472 => x"30",
         15473 => x"25",
         15474 => x"00",
         15475 => x"44",
         15476 => x"30",
         15477 => x"25",
         15478 => x"00",
         15479 => x"48",
         15480 => x"30",
         15481 => x"00",
         15482 => x"4e",
         15483 => x"65",
         15484 => x"64",
         15485 => x"6e",
         15486 => x"00",
         15487 => x"53",
         15488 => x"22",
         15489 => x"3e",
         15490 => x"00",
         15491 => x"2b",
         15492 => x"5b",
         15493 => x"46",
         15494 => x"46",
         15495 => x"32",
         15496 => x"eb",
         15497 => x"53",
         15498 => x"35",
         15499 => x"4e",
         15500 => x"41",
         15501 => x"20",
         15502 => x"41",
         15503 => x"20",
         15504 => x"4e",
         15505 => x"41",
         15506 => x"20",
         15507 => x"41",
         15508 => x"20",
         15509 => x"00",
         15510 => x"00",
         15511 => x"00",
         15512 => x"00",
         15513 => x"01",
         15514 => x"09",
         15515 => x"14",
         15516 => x"1e",
         15517 => x"80",
         15518 => x"8e",
         15519 => x"45",
         15520 => x"49",
         15521 => x"90",
         15522 => x"99",
         15523 => x"59",
         15524 => x"9c",
         15525 => x"41",
         15526 => x"a5",
         15527 => x"a8",
         15528 => x"ac",
         15529 => x"b0",
         15530 => x"b4",
         15531 => x"b8",
         15532 => x"bc",
         15533 => x"c0",
         15534 => x"c4",
         15535 => x"c8",
         15536 => x"cc",
         15537 => x"d0",
         15538 => x"d4",
         15539 => x"d8",
         15540 => x"dc",
         15541 => x"e0",
         15542 => x"e4",
         15543 => x"e8",
         15544 => x"ec",
         15545 => x"f0",
         15546 => x"f4",
         15547 => x"f8",
         15548 => x"fc",
         15549 => x"2b",
         15550 => x"3d",
         15551 => x"5c",
         15552 => x"3c",
         15553 => x"7f",
         15554 => x"00",
         15555 => x"00",
         15556 => x"01",
         15557 => x"00",
         15558 => x"00",
         15559 => x"00",
         15560 => x"00",
         15561 => x"00",
         15562 => x"00",
         15563 => x"00",
         15564 => x"00",
         15565 => x"00",
         15566 => x"00",
         15567 => x"00",
         15568 => x"00",
         15569 => x"00",
         15570 => x"00",
         15571 => x"00",
         15572 => x"00",
         15573 => x"00",
         15574 => x"00",
         15575 => x"00",
         15576 => x"00",
         15577 => x"20",
         15578 => x"00",
         15579 => x"00",
         15580 => x"00",
         15581 => x"00",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"00",
         15586 => x"25",
         15587 => x"25",
         15588 => x"25",
         15589 => x"25",
         15590 => x"25",
         15591 => x"25",
         15592 => x"25",
         15593 => x"25",
         15594 => x"25",
         15595 => x"25",
         15596 => x"25",
         15597 => x"25",
         15598 => x"25",
         15599 => x"25",
         15600 => x"25",
         15601 => x"25",
         15602 => x"25",
         15603 => x"25",
         15604 => x"25",
         15605 => x"25",
         15606 => x"25",
         15607 => x"25",
         15608 => x"25",
         15609 => x"25",
         15610 => x"03",
         15611 => x"03",
         15612 => x"03",
         15613 => x"00",
         15614 => x"03",
         15615 => x"03",
         15616 => x"22",
         15617 => x"03",
         15618 => x"22",
         15619 => x"22",
         15620 => x"23",
         15621 => x"00",
         15622 => x"00",
         15623 => x"00",
         15624 => x"20",
         15625 => x"25",
         15626 => x"00",
         15627 => x"00",
         15628 => x"00",
         15629 => x"00",
         15630 => x"01",
         15631 => x"01",
         15632 => x"01",
         15633 => x"01",
         15634 => x"01",
         15635 => x"01",
         15636 => x"00",
         15637 => x"01",
         15638 => x"01",
         15639 => x"01",
         15640 => x"01",
         15641 => x"01",
         15642 => x"01",
         15643 => x"01",
         15644 => x"01",
         15645 => x"01",
         15646 => x"01",
         15647 => x"01",
         15648 => x"01",
         15649 => x"01",
         15650 => x"01",
         15651 => x"01",
         15652 => x"01",
         15653 => x"01",
         15654 => x"01",
         15655 => x"01",
         15656 => x"01",
         15657 => x"01",
         15658 => x"01",
         15659 => x"01",
         15660 => x"01",
         15661 => x"01",
         15662 => x"01",
         15663 => x"01",
         15664 => x"01",
         15665 => x"01",
         15666 => x"01",
         15667 => x"01",
         15668 => x"01",
         15669 => x"01",
         15670 => x"01",
         15671 => x"01",
         15672 => x"01",
         15673 => x"01",
         15674 => x"01",
         15675 => x"01",
         15676 => x"01",
         15677 => x"01",
         15678 => x"01",
         15679 => x"00",
         15680 => x"01",
         15681 => x"01",
         15682 => x"02",
         15683 => x"02",
         15684 => x"2c",
         15685 => x"02",
         15686 => x"2c",
         15687 => x"02",
         15688 => x"02",
         15689 => x"01",
         15690 => x"00",
         15691 => x"01",
         15692 => x"01",
         15693 => x"02",
         15694 => x"02",
         15695 => x"02",
         15696 => x"02",
         15697 => x"01",
         15698 => x"02",
         15699 => x"02",
         15700 => x"02",
         15701 => x"01",
         15702 => x"02",
         15703 => x"02",
         15704 => x"02",
         15705 => x"02",
         15706 => x"01",
         15707 => x"02",
         15708 => x"02",
         15709 => x"02",
         15710 => x"02",
         15711 => x"02",
         15712 => x"02",
         15713 => x"01",
         15714 => x"02",
         15715 => x"02",
         15716 => x"02",
         15717 => x"01",
         15718 => x"01",
         15719 => x"02",
         15720 => x"02",
         15721 => x"02",
         15722 => x"01",
         15723 => x"00",
         15724 => x"03",
         15725 => x"03",
         15726 => x"03",
         15727 => x"03",
         15728 => x"03",
         15729 => x"03",
         15730 => x"03",
         15731 => x"03",
         15732 => x"03",
         15733 => x"03",
         15734 => x"03",
         15735 => x"01",
         15736 => x"00",
         15737 => x"03",
         15738 => x"03",
         15739 => x"03",
         15740 => x"03",
         15741 => x"03",
         15742 => x"03",
         15743 => x"07",
         15744 => x"01",
         15745 => x"01",
         15746 => x"01",
         15747 => x"00",
         15748 => x"04",
         15749 => x"05",
         15750 => x"00",
         15751 => x"1d",
         15752 => x"2c",
         15753 => x"01",
         15754 => x"01",
         15755 => x"06",
         15756 => x"06",
         15757 => x"06",
         15758 => x"06",
         15759 => x"06",
         15760 => x"00",
         15761 => x"1f",
         15762 => x"1f",
         15763 => x"1f",
         15764 => x"1f",
         15765 => x"1f",
         15766 => x"1f",
         15767 => x"1f",
         15768 => x"1f",
         15769 => x"1f",
         15770 => x"1f",
         15771 => x"1f",
         15772 => x"1f",
         15773 => x"1f",
         15774 => x"1f",
         15775 => x"1f",
         15776 => x"1f",
         15777 => x"1f",
         15778 => x"1f",
         15779 => x"1f",
         15780 => x"1f",
         15781 => x"06",
         15782 => x"06",
         15783 => x"00",
         15784 => x"1f",
         15785 => x"1f",
         15786 => x"00",
         15787 => x"21",
         15788 => x"21",
         15789 => x"21",
         15790 => x"05",
         15791 => x"04",
         15792 => x"01",
         15793 => x"01",
         15794 => x"01",
         15795 => x"01",
         15796 => x"08",
         15797 => x"03",
         15798 => x"00",
         15799 => x"00",
         15800 => x"01",
         15801 => x"00",
         15802 => x"00",
         15803 => x"00",
         15804 => x"01",
         15805 => x"00",
         15806 => x"00",
         15807 => x"00",
         15808 => x"01",
         15809 => x"00",
         15810 => x"00",
         15811 => x"00",
         15812 => x"01",
         15813 => x"00",
         15814 => x"00",
         15815 => x"00",
         15816 => x"01",
         15817 => x"00",
         15818 => x"00",
         15819 => x"00",
         15820 => x"01",
         15821 => x"00",
         15822 => x"00",
         15823 => x"00",
         15824 => x"01",
         15825 => x"00",
         15826 => x"00",
         15827 => x"00",
         15828 => x"01",
         15829 => x"00",
         15830 => x"00",
         15831 => x"00",
         15832 => x"01",
         15833 => x"00",
         15834 => x"00",
         15835 => x"00",
         15836 => x"01",
         15837 => x"00",
         15838 => x"00",
         15839 => x"00",
         15840 => x"01",
         15841 => x"00",
         15842 => x"00",
         15843 => x"00",
         15844 => x"01",
         15845 => x"00",
         15846 => x"00",
         15847 => x"00",
         15848 => x"01",
         15849 => x"00",
         15850 => x"00",
         15851 => x"00",
         15852 => x"01",
         15853 => x"00",
         15854 => x"00",
         15855 => x"00",
         15856 => x"01",
         15857 => x"00",
         15858 => x"00",
         15859 => x"00",
         15860 => x"01",
         15861 => x"00",
         15862 => x"00",
         15863 => x"00",
         15864 => x"01",
         15865 => x"00",
         15866 => x"00",
         15867 => x"00",
         15868 => x"01",
         15869 => x"00",
         15870 => x"00",
         15871 => x"00",
         15872 => x"01",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"01",
         15877 => x"00",
         15878 => x"00",
         15879 => x"00",
         15880 => x"01",
         15881 => x"00",
         15882 => x"00",
         15883 => x"00",
         15884 => x"01",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"01",
         15889 => x"00",
         15890 => x"00",
         15891 => x"00",
         15892 => x"01",
         15893 => x"00",
         15894 => x"00",
         15895 => x"00",
         15896 => x"01",
         15897 => x"00",
         15898 => x"00",
         15899 => x"00",
         15900 => x"01",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"01",
         15905 => x"00",
         15906 => x"00",
         15907 => x"00",
         15908 => x"01",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"00",
         15913 => x"00",
         15914 => x"00",
         15915 => x"00",
         15916 => x"00",
         15917 => x"00",
         15918 => x"00",
         15919 => x"00",
         15920 => x"01",
         15921 => x"01",
         15922 => x"00",
         15923 => x"00",
         15924 => x"00",
         15925 => x"00",
         15926 => x"05",
         15927 => x"05",
         15928 => x"05",
         15929 => x"00",
         15930 => x"01",
         15931 => x"01",
         15932 => x"01",
         15933 => x"01",
         15934 => x"00",
         15935 => x"00",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"00",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"00",
         15957 => x"00",
         15958 => x"00",
         15959 => x"01",
         15960 => x"00",
         15961 => x"01",
         15962 => x"00",
         15963 => x"02",
         15964 => x"00",
         15965 => x"1b",
         15966 => x"f0",
         15967 => x"79",
         15968 => x"5d",
         15969 => x"71",
         15970 => x"75",
         15971 => x"69",
         15972 => x"6d",
         15973 => x"61",
         15974 => x"65",
         15975 => x"31",
         15976 => x"35",
         15977 => x"5c",
         15978 => x"30",
         15979 => x"f6",
         15980 => x"f1",
         15981 => x"08",
         15982 => x"f0",
         15983 => x"80",
         15984 => x"84",
         15985 => x"1b",
         15986 => x"f0",
         15987 => x"59",
         15988 => x"5d",
         15989 => x"51",
         15990 => x"55",
         15991 => x"49",
         15992 => x"4d",
         15993 => x"41",
         15994 => x"45",
         15995 => x"31",
         15996 => x"35",
         15997 => x"5c",
         15998 => x"30",
         15999 => x"f6",
         16000 => x"f1",
         16001 => x"08",
         16002 => x"f0",
         16003 => x"80",
         16004 => x"84",
         16005 => x"1b",
         16006 => x"f0",
         16007 => x"59",
         16008 => x"7d",
         16009 => x"51",
         16010 => x"55",
         16011 => x"49",
         16012 => x"4d",
         16013 => x"41",
         16014 => x"45",
         16015 => x"21",
         16016 => x"25",
         16017 => x"7c",
         16018 => x"20",
         16019 => x"f7",
         16020 => x"f9",
         16021 => x"fb",
         16022 => x"f0",
         16023 => x"85",
         16024 => x"89",
         16025 => x"1b",
         16026 => x"f0",
         16027 => x"19",
         16028 => x"1d",
         16029 => x"11",
         16030 => x"15",
         16031 => x"09",
         16032 => x"0d",
         16033 => x"01",
         16034 => x"05",
         16035 => x"f0",
         16036 => x"f0",
         16037 => x"f0",
         16038 => x"f0",
         16039 => x"f0",
         16040 => x"f0",
         16041 => x"f0",
         16042 => x"f0",
         16043 => x"80",
         16044 => x"84",
         16045 => x"bf",
         16046 => x"f0",
         16047 => x"35",
         16048 => x"b7",
         16049 => x"7c",
         16050 => x"39",
         16051 => x"3d",
         16052 => x"1d",
         16053 => x"46",
         16054 => x"74",
         16055 => x"3f",
         16056 => x"7a",
         16057 => x"d3",
         16058 => x"9d",
         16059 => x"c6",
         16060 => x"c3",
         16061 => x"f0",
         16062 => x"f0",
         16063 => x"80",
         16064 => x"84",
         16065 => x"00",
         16066 => x"00",
         16067 => x"00",
         16068 => x"00",
         16069 => x"00",
         16070 => x"00",
         16071 => x"00",
         16072 => x"00",
         16073 => x"00",
         16074 => x"00",
         16075 => x"00",
         16076 => x"00",
         16077 => x"00",
         16078 => x"00",
         16079 => x"00",
         16080 => x"00",
         16081 => x"00",
         16082 => x"00",
         16083 => x"00",
         16084 => x"00",
         16085 => x"00",
         16086 => x"00",
         16087 => x"00",
         16088 => x"00",
         16089 => x"00",
         16090 => x"00",
         16091 => x"00",
         16092 => x"f8",
         16093 => x"00",
         16094 => x"f3",
         16095 => x"00",
         16096 => x"f4",
         16097 => x"00",
         16098 => x"f1",
         16099 => x"00",
         16100 => x"f2",
         16101 => x"00",
         16102 => x"80",
         16103 => x"00",
         16104 => x"81",
         16105 => x"00",
         16106 => x"82",
         16107 => x"00",
         16108 => x"83",
         16109 => x"00",
         16110 => x"84",
         16111 => x"00",
         16112 => x"85",
         16113 => x"00",
         16114 => x"86",
         16115 => x"00",
         16116 => x"87",
         16117 => x"00",
         16118 => x"88",
         16119 => x"00",
         16120 => x"89",
         16121 => x"00",
         16122 => x"f6",
         16123 => x"00",
         16124 => x"7f",
         16125 => x"00",
         16126 => x"f9",
         16127 => x"00",
         16128 => x"e0",
         16129 => x"00",
         16130 => x"e1",
         16131 => x"00",
         16132 => x"71",
         16133 => x"00",
         16134 => x"00",
         16135 => x"00",
         16136 => x"00",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"50",
         18135 => x"00",
         18136 => x"cc",
         18137 => x"ce",
         18138 => x"f8",
         18139 => x"fc",
         18140 => x"e1",
         18141 => x"c4",
         18142 => x"e3",
         18143 => x"eb",
         18144 => x"00",
         18145 => x"64",
         18146 => x"68",
         18147 => x"2f",
         18148 => x"20",
         18149 => x"24",
         18150 => x"28",
         18151 => x"51",
         18152 => x"55",
         18153 => x"04",
         18154 => x"08",
         18155 => x"0c",
         18156 => x"10",
         18157 => x"14",
         18158 => x"18",
         18159 => x"59",
         18160 => x"c7",
         18161 => x"84",
         18162 => x"88",
         18163 => x"8c",
         18164 => x"90",
         18165 => x"94",
         18166 => x"98",
         18167 => x"80",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
