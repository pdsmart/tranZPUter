-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"ac",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c5",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c7",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"e4",
           386 => x"d4",
           387 => x"e4",
           388 => x"90",
           389 => x"e4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"84",
           396 => x"82",
           397 => x"af",
           398 => x"d6",
           399 => x"80",
           400 => x"d6",
           401 => x"ad",
           402 => x"e4",
           403 => x"90",
           404 => x"e4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"84",
           419 => x"82",
           420 => x"96",
           421 => x"d6",
           422 => x"80",
           423 => x"d6",
           424 => x"cd",
           425 => x"e4",
           426 => x"90",
           427 => x"e4",
           428 => x"fa",
           429 => x"e4",
           430 => x"90",
           431 => x"e4",
           432 => x"c9",
           433 => x"e4",
           434 => x"90",
           435 => x"e4",
           436 => x"99",
           437 => x"e4",
           438 => x"90",
           439 => x"e4",
           440 => x"90",
           441 => x"e4",
           442 => x"90",
           443 => x"e4",
           444 => x"c3",
           445 => x"e4",
           446 => x"90",
           447 => x"e4",
           448 => x"ad",
           449 => x"e4",
           450 => x"90",
           451 => x"e4",
           452 => x"ac",
           453 => x"e4",
           454 => x"90",
           455 => x"e4",
           456 => x"92",
           457 => x"e4",
           458 => x"90",
           459 => x"e4",
           460 => x"92",
           461 => x"e4",
           462 => x"90",
           463 => x"e4",
           464 => x"ea",
           465 => x"e4",
           466 => x"90",
           467 => x"e4",
           468 => x"d3",
           469 => x"e4",
           470 => x"90",
           471 => x"e4",
           472 => x"89",
           473 => x"e4",
           474 => x"90",
           475 => x"e4",
           476 => x"8d",
           477 => x"e4",
           478 => x"90",
           479 => x"e4",
           480 => x"ad",
           481 => x"e4",
           482 => x"90",
           483 => x"e4",
           484 => x"cc",
           485 => x"e4",
           486 => x"90",
           487 => x"e4",
           488 => x"c0",
           489 => x"e4",
           490 => x"90",
           491 => x"e4",
           492 => x"a2",
           493 => x"e4",
           494 => x"90",
           495 => x"e4",
           496 => x"9c",
           497 => x"e4",
           498 => x"90",
           499 => x"e4",
           500 => x"d2",
           501 => x"e4",
           502 => x"90",
           503 => x"e4",
           504 => x"a1",
           505 => x"e4",
           506 => x"90",
           507 => x"e4",
           508 => x"a2",
           509 => x"e4",
           510 => x"90",
           511 => x"e4",
           512 => x"8c",
           513 => x"e4",
           514 => x"90",
           515 => x"e4",
           516 => x"e5",
           517 => x"e4",
           518 => x"90",
           519 => x"e4",
           520 => x"90",
           521 => x"e4",
           522 => x"90",
           523 => x"e4",
           524 => x"a9",
           525 => x"e4",
           526 => x"90",
           527 => x"e4",
           528 => x"93",
           529 => x"e4",
           530 => x"90",
           531 => x"e4",
           532 => x"9e",
           533 => x"e4",
           534 => x"90",
           535 => x"e4",
           536 => x"a5",
           537 => x"e4",
           538 => x"90",
           539 => x"e4",
           540 => x"cc",
           541 => x"e4",
           542 => x"90",
           543 => x"e4",
           544 => x"91",
           545 => x"e4",
           546 => x"90",
           547 => x"e4",
           548 => x"c6",
           549 => x"e4",
           550 => x"90",
           551 => x"e4",
           552 => x"b2",
           553 => x"e4",
           554 => x"90",
           555 => x"e4",
           556 => x"d4",
           557 => x"e4",
           558 => x"90",
           559 => x"e4",
           560 => x"be",
           561 => x"e4",
           562 => x"90",
           563 => x"e4",
           564 => x"a2",
           565 => x"e4",
           566 => x"90",
           567 => x"e4",
           568 => x"c2",
           569 => x"e4",
           570 => x"90",
           571 => x"e4",
           572 => x"e6",
           573 => x"e4",
           574 => x"90",
           575 => x"e4",
           576 => x"c9",
           577 => x"e4",
           578 => x"90",
           579 => x"e4",
           580 => x"bf",
           581 => x"e4",
           582 => x"90",
           583 => x"e4",
           584 => x"e8",
           585 => x"e4",
           586 => x"90",
           587 => x"e4",
           588 => x"90",
           589 => x"e4",
           590 => x"90",
           591 => x"e4",
           592 => x"88",
           593 => x"e4",
           594 => x"90",
           595 => x"e4",
           596 => x"d2",
           597 => x"e4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"d8",
           623 => x"c4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"e4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"d6",
           637 => x"05",
           638 => x"d6",
           639 => x"05",
           640 => x"f2",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"e4",
           652 => x"d6",
           653 => x"3d",
           654 => x"e4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"d6",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"d6",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"d6",
           675 => x"05",
           676 => x"e4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"d6",
           683 => x"05",
           684 => x"90",
           685 => x"d8",
           686 => x"d6",
           687 => x"05",
           688 => x"d6",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"d6",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"d6",
           709 => x"05",
           710 => x"72",
           711 => x"e4",
           712 => x"08",
           713 => x"e4",
           714 => x"0c",
           715 => x"e4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"e4",
           722 => x"0d",
           723 => x"d6",
           724 => x"05",
           725 => x"e4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"d6",
           730 => x"05",
           731 => x"e4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"e4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"e4",
           756 => x"d6",
           757 => x"3d",
           758 => x"e4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"d6",
           769 => x"82",
           770 => x"f8",
           771 => x"d6",
           772 => x"05",
           773 => x"d6",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"e4",
           779 => x"0d",
           780 => x"d6",
           781 => x"05",
           782 => x"e4",
           783 => x"08",
           784 => x"8c",
           785 => x"d6",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"e4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"e4",
           804 => x"08",
           805 => x"d6",
           806 => x"05",
           807 => x"e4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"e4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"d6",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"e4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"d6",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"d6",
           863 => x"05",
           864 => x"e4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"e4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"d6",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"e4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"d6",
           889 => x"05",
           890 => x"e4",
           891 => x"33",
           892 => x"d6",
           893 => x"05",
           894 => x"d6",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"bc",
           901 => x"51",
           902 => x"72",
           903 => x"e4",
           904 => x"22",
           905 => x"51",
           906 => x"d6",
           907 => x"05",
           908 => x"e4",
           909 => x"22",
           910 => x"51",
           911 => x"d6",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"d6",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"d6",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"e4",
           930 => x"23",
           931 => x"d6",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"e4",
           938 => x"23",
           939 => x"bf",
           940 => x"e4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"d6",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"e4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"e4",
           969 => x"0c",
           970 => x"d6",
           971 => x"05",
           972 => x"e4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"d6",
           982 => x"05",
           983 => x"a4",
           984 => x"d6",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"e4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"d6",
           993 => x"05",
           994 => x"e4",
           995 => x"22",
           996 => x"e4",
           997 => x"22",
           998 => x"54",
           999 => x"d6",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"e4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"d6",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"e4",
          1020 => x"08",
          1021 => x"ec",
          1022 => x"d8",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"e4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"e4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"e4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"d6",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"d6",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"e4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"d6",
          1072 => x"05",
          1073 => x"e4",
          1074 => x"08",
          1075 => x"e4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"d6",
          1081 => x"05",
          1082 => x"39",
          1083 => x"d6",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"e4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"e4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"d6",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"d6",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"d6",
          1127 => x"d6",
          1128 => x"05",
          1129 => x"e4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"d6",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"d6",
          1147 => x"05",
          1148 => x"33",
          1149 => x"e4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"e4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"e4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"e4",
          1172 => x"08",
          1173 => x"d6",
          1174 => x"d8",
          1175 => x"d6",
          1176 => x"05",
          1177 => x"d6",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"e4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"e4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"e4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"d6",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"d6",
          1225 => x"05",
          1226 => x"e4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"d6",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"e4",
          1247 => x"33",
          1248 => x"e4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"d6",
          1252 => x"05",
          1253 => x"e4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"d6",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"e4",
          1269 => x"23",
          1270 => x"d6",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"e4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"e4",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"e4",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"d6",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"d6",
          1381 => x"05",
          1382 => x"54",
          1383 => x"d6",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"d6",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"e4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"d6",
          1397 => x"05",
          1398 => x"d6",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"d6",
          1407 => x"05",
          1408 => x"51",
          1409 => x"d6",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"e4",
          1420 => x"08",
          1421 => x"d6",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"d6",
          1430 => x"05",
          1431 => x"51",
          1432 => x"d6",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"e4",
          1444 => x"08",
          1445 => x"d6",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"e4",
          1452 => x"08",
          1453 => x"e4",
          1454 => x"08",
          1455 => x"d6",
          1456 => x"05",
          1457 => x"e4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"e4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"d6",
          1479 => x"05",
          1480 => x"d6",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"e4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"e4",
          1496 => x"34",
          1497 => x"d6",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"d6",
          1506 => x"05",
          1507 => x"08",
          1508 => x"e4",
          1509 => x"0c",
          1510 => x"d6",
          1511 => x"05",
          1512 => x"d8",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"e4",
          1516 => x"d6",
          1517 => x"3d",
          1518 => x"b8",
          1519 => x"d6",
          1520 => x"05",
          1521 => x"d6",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"d8",
          1525 => x"d6",
          1526 => x"85",
          1527 => x"d6",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"e4",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"d6",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"e4",
          1549 => x"0c",
          1550 => x"d6",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"f2",
          1567 => x"f2",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"d6",
          1582 => x"3d",
          1583 => x"e4",
          1584 => x"d6",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"d6",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"d6",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"e4",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"d6",
          1625 => x"05",
          1626 => x"d6",
          1627 => x"05",
          1628 => x"d6",
          1629 => x"05",
          1630 => x"d8",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"e4",
          1634 => x"d6",
          1635 => x"3d",
          1636 => x"bc",
          1637 => x"d6",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"d8",
          1642 => x"3d",
          1643 => x"e4",
          1644 => x"d6",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"d6",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"e4",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"e4",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"d6",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"d6",
          1689 => x"05",
          1690 => x"d6",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"d6",
          1696 => x"72",
          1697 => x"d6",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"e4",
          1702 => x"08",
          1703 => x"e4",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"d6",
          1707 => x"05",
          1708 => x"e4",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"e4",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"e4",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"d6",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"d6",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"e4",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"e4",
          1761 => x"08",
          1762 => x"d6",
          1763 => x"05",
          1764 => x"e4",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"d6",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"d6",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"d8",
          1783 => x"d6",
          1784 => x"05",
          1785 => x"d6",
          1786 => x"05",
          1787 => x"80",
          1788 => x"d6",
          1789 => x"05",
          1790 => x"e4",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"d6",
          1795 => x"05",
          1796 => x"d6",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"d6",
          1810 => x"05",
          1811 => x"d6",
          1812 => x"05",
          1813 => x"34",
          1814 => x"d6",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"d6",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"d6",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"d6",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"d6",
          1836 => x"05",
          1837 => x"e4",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"d6",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"e4",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"e4",
          1853 => x"08",
          1854 => x"90",
          1855 => x"e4",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"d6",
          1863 => x"05",
          1864 => x"d6",
          1865 => x"05",
          1866 => x"e4",
          1867 => x"08",
          1868 => x"d6",
          1869 => x"05",
          1870 => x"e4",
          1871 => x"08",
          1872 => x"d6",
          1873 => x"05",
          1874 => x"e4",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"e4",
          1878 => x"08",
          1879 => x"d6",
          1880 => x"05",
          1881 => x"e4",
          1882 => x"08",
          1883 => x"d6",
          1884 => x"05",
          1885 => x"e4",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"e4",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"e4",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"e4",
          1905 => x"08",
          1906 => x"d6",
          1907 => x"05",
          1908 => x"e4",
          1909 => x"08",
          1910 => x"71",
          1911 => x"e4",
          1912 => x"08",
          1913 => x"d6",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"e4",
          1922 => x"d6",
          1923 => x"3d",
          1924 => x"e4",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"e4",
          1931 => x"08",
          1932 => x"d6",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"d6",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"d6",
          1942 => x"05",
          1943 => x"e4",
          1944 => x"08",
          1945 => x"d6",
          1946 => x"84",
          1947 => x"d6",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"d6",
          1954 => x"05",
          1955 => x"e4",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"e4",
          1978 => x"d6",
          1979 => x"3d",
          1980 => x"e4",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"d6",
          1986 => x"05",
          1987 => x"e4",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"e4",
          1991 => x"08",
          1992 => x"d6",
          1993 => x"05",
          1994 => x"e4",
          1995 => x"08",
          1996 => x"d6",
          1997 => x"05",
          1998 => x"e4",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"d6",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"d6",
          2008 => x"05",
          2009 => x"71",
          2010 => x"d6",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"e4",
          2016 => x"08",
          2017 => x"d8",
          2018 => x"3d",
          2019 => x"e4",
          2020 => x"d6",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"d6",
          2024 => x"05",
          2025 => x"81",
          2026 => x"d6",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"e4",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"e4",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"d6",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"e4",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"d6",
          2059 => x"05",
          2060 => x"80",
          2061 => x"d6",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"d6",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"e4",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"e4",
          2079 => x"08",
          2080 => x"d6",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"d6",
          2090 => x"05",
          2091 => x"d8",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"e4",
          2095 => x"d6",
          2096 => x"3d",
          2097 => x"e4",
          2098 => x"08",
          2099 => x"e4",
          2100 => x"08",
          2101 => x"3f",
          2102 => x"08",
          2103 => x"e4",
          2104 => x"0c",
          2105 => x"08",
          2106 => x"81",
          2107 => x"51",
          2108 => x"f4",
          2109 => x"d8",
          2110 => x"d6",
          2111 => x"05",
          2112 => x"d6",
          2113 => x"05",
          2114 => x"80",
          2115 => x"e4",
          2116 => x"0c",
          2117 => x"d6",
          2118 => x"05",
          2119 => x"e4",
          2120 => x"08",
          2121 => x"74",
          2122 => x"e4",
          2123 => x"08",
          2124 => x"e4",
          2125 => x"08",
          2126 => x"e4",
          2127 => x"08",
          2128 => x"3f",
          2129 => x"08",
          2130 => x"e4",
          2131 => x"0c",
          2132 => x"e4",
          2133 => x"08",
          2134 => x"0c",
          2135 => x"82",
          2136 => x"04",
          2137 => x"08",
          2138 => x"e4",
          2139 => x"0d",
          2140 => x"08",
          2141 => x"82",
          2142 => x"f8",
          2143 => x"d6",
          2144 => x"05",
          2145 => x"80",
          2146 => x"e4",
          2147 => x"0c",
          2148 => x"82",
          2149 => x"f8",
          2150 => x"71",
          2151 => x"e4",
          2152 => x"08",
          2153 => x"d6",
          2154 => x"05",
          2155 => x"ff",
          2156 => x"70",
          2157 => x"38",
          2158 => x"08",
          2159 => x"ff",
          2160 => x"e4",
          2161 => x"0c",
          2162 => x"08",
          2163 => x"ff",
          2164 => x"ff",
          2165 => x"d6",
          2166 => x"05",
          2167 => x"82",
          2168 => x"f8",
          2169 => x"d6",
          2170 => x"05",
          2171 => x"e4",
          2172 => x"08",
          2173 => x"d6",
          2174 => x"05",
          2175 => x"d6",
          2176 => x"05",
          2177 => x"d8",
          2178 => x"0d",
          2179 => x"0c",
          2180 => x"e4",
          2181 => x"d6",
          2182 => x"3d",
          2183 => x"e4",
          2184 => x"08",
          2185 => x"08",
          2186 => x"82",
          2187 => x"90",
          2188 => x"2e",
          2189 => x"82",
          2190 => x"90",
          2191 => x"05",
          2192 => x"08",
          2193 => x"82",
          2194 => x"90",
          2195 => x"05",
          2196 => x"08",
          2197 => x"82",
          2198 => x"90",
          2199 => x"2e",
          2200 => x"d6",
          2201 => x"05",
          2202 => x"82",
          2203 => x"fc",
          2204 => x"52",
          2205 => x"82",
          2206 => x"fc",
          2207 => x"05",
          2208 => x"08",
          2209 => x"ff",
          2210 => x"d6",
          2211 => x"05",
          2212 => x"d6",
          2213 => x"84",
          2214 => x"d6",
          2215 => x"82",
          2216 => x"02",
          2217 => x"0c",
          2218 => x"80",
          2219 => x"e4",
          2220 => x"0c",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"88",
          2225 => x"82",
          2226 => x"88",
          2227 => x"0b",
          2228 => x"08",
          2229 => x"82",
          2230 => x"fc",
          2231 => x"38",
          2232 => x"d6",
          2233 => x"05",
          2234 => x"e4",
          2235 => x"08",
          2236 => x"08",
          2237 => x"82",
          2238 => x"8c",
          2239 => x"25",
          2240 => x"d6",
          2241 => x"05",
          2242 => x"d6",
          2243 => x"05",
          2244 => x"82",
          2245 => x"f0",
          2246 => x"d6",
          2247 => x"05",
          2248 => x"81",
          2249 => x"e4",
          2250 => x"0c",
          2251 => x"08",
          2252 => x"82",
          2253 => x"fc",
          2254 => x"53",
          2255 => x"08",
          2256 => x"52",
          2257 => x"08",
          2258 => x"51",
          2259 => x"82",
          2260 => x"70",
          2261 => x"08",
          2262 => x"54",
          2263 => x"08",
          2264 => x"80",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"d6",
          2270 => x"05",
          2271 => x"d6",
          2272 => x"89",
          2273 => x"d6",
          2274 => x"82",
          2275 => x"02",
          2276 => x"0c",
          2277 => x"80",
          2278 => x"e4",
          2279 => x"0c",
          2280 => x"08",
          2281 => x"80",
          2282 => x"82",
          2283 => x"88",
          2284 => x"82",
          2285 => x"88",
          2286 => x"0b",
          2287 => x"08",
          2288 => x"82",
          2289 => x"8c",
          2290 => x"25",
          2291 => x"d6",
          2292 => x"05",
          2293 => x"d6",
          2294 => x"05",
          2295 => x"82",
          2296 => x"8c",
          2297 => x"82",
          2298 => x"88",
          2299 => x"81",
          2300 => x"d6",
          2301 => x"82",
          2302 => x"f8",
          2303 => x"82",
          2304 => x"fc",
          2305 => x"2e",
          2306 => x"d6",
          2307 => x"05",
          2308 => x"d6",
          2309 => x"05",
          2310 => x"e4",
          2311 => x"08",
          2312 => x"d8",
          2313 => x"3d",
          2314 => x"e4",
          2315 => x"d6",
          2316 => x"82",
          2317 => x"fd",
          2318 => x"53",
          2319 => x"08",
          2320 => x"52",
          2321 => x"08",
          2322 => x"51",
          2323 => x"82",
          2324 => x"70",
          2325 => x"0c",
          2326 => x"0d",
          2327 => x"0c",
          2328 => x"e4",
          2329 => x"d6",
          2330 => x"3d",
          2331 => x"82",
          2332 => x"8c",
          2333 => x"82",
          2334 => x"88",
          2335 => x"93",
          2336 => x"d8",
          2337 => x"d6",
          2338 => x"85",
          2339 => x"d6",
          2340 => x"82",
          2341 => x"02",
          2342 => x"0c",
          2343 => x"81",
          2344 => x"e4",
          2345 => x"0c",
          2346 => x"d6",
          2347 => x"05",
          2348 => x"e4",
          2349 => x"08",
          2350 => x"08",
          2351 => x"27",
          2352 => x"d6",
          2353 => x"05",
          2354 => x"ae",
          2355 => x"82",
          2356 => x"8c",
          2357 => x"a2",
          2358 => x"e4",
          2359 => x"08",
          2360 => x"e4",
          2361 => x"0c",
          2362 => x"08",
          2363 => x"10",
          2364 => x"08",
          2365 => x"ff",
          2366 => x"d6",
          2367 => x"05",
          2368 => x"80",
          2369 => x"d6",
          2370 => x"05",
          2371 => x"e4",
          2372 => x"08",
          2373 => x"82",
          2374 => x"88",
          2375 => x"d6",
          2376 => x"05",
          2377 => x"d6",
          2378 => x"05",
          2379 => x"e4",
          2380 => x"08",
          2381 => x"08",
          2382 => x"07",
          2383 => x"08",
          2384 => x"82",
          2385 => x"fc",
          2386 => x"2a",
          2387 => x"08",
          2388 => x"82",
          2389 => x"8c",
          2390 => x"2a",
          2391 => x"08",
          2392 => x"ff",
          2393 => x"d6",
          2394 => x"05",
          2395 => x"93",
          2396 => x"e4",
          2397 => x"08",
          2398 => x"e4",
          2399 => x"0c",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"82",
          2403 => x"f4",
          2404 => x"82",
          2405 => x"f4",
          2406 => x"d6",
          2407 => x"3d",
          2408 => x"e4",
          2409 => x"d6",
          2410 => x"82",
          2411 => x"f7",
          2412 => x"0b",
          2413 => x"08",
          2414 => x"82",
          2415 => x"8c",
          2416 => x"80",
          2417 => x"d6",
          2418 => x"05",
          2419 => x"51",
          2420 => x"53",
          2421 => x"e4",
          2422 => x"34",
          2423 => x"06",
          2424 => x"2e",
          2425 => x"91",
          2426 => x"e4",
          2427 => x"08",
          2428 => x"05",
          2429 => x"ce",
          2430 => x"e4",
          2431 => x"33",
          2432 => x"2e",
          2433 => x"a4",
          2434 => x"82",
          2435 => x"f0",
          2436 => x"d6",
          2437 => x"05",
          2438 => x"81",
          2439 => x"70",
          2440 => x"72",
          2441 => x"e4",
          2442 => x"34",
          2443 => x"08",
          2444 => x"53",
          2445 => x"09",
          2446 => x"dc",
          2447 => x"e4",
          2448 => x"08",
          2449 => x"05",
          2450 => x"08",
          2451 => x"33",
          2452 => x"08",
          2453 => x"82",
          2454 => x"f8",
          2455 => x"d6",
          2456 => x"05",
          2457 => x"e4",
          2458 => x"08",
          2459 => x"b6",
          2460 => x"e4",
          2461 => x"08",
          2462 => x"84",
          2463 => x"39",
          2464 => x"d6",
          2465 => x"05",
          2466 => x"e4",
          2467 => x"08",
          2468 => x"05",
          2469 => x"08",
          2470 => x"33",
          2471 => x"08",
          2472 => x"81",
          2473 => x"0b",
          2474 => x"08",
          2475 => x"82",
          2476 => x"88",
          2477 => x"08",
          2478 => x"0c",
          2479 => x"53",
          2480 => x"d6",
          2481 => x"05",
          2482 => x"39",
          2483 => x"08",
          2484 => x"53",
          2485 => x"8d",
          2486 => x"82",
          2487 => x"ec",
          2488 => x"80",
          2489 => x"e4",
          2490 => x"33",
          2491 => x"27",
          2492 => x"d6",
          2493 => x"05",
          2494 => x"b9",
          2495 => x"8d",
          2496 => x"82",
          2497 => x"ec",
          2498 => x"d8",
          2499 => x"82",
          2500 => x"f4",
          2501 => x"39",
          2502 => x"08",
          2503 => x"53",
          2504 => x"90",
          2505 => x"e4",
          2506 => x"33",
          2507 => x"26",
          2508 => x"39",
          2509 => x"d6",
          2510 => x"05",
          2511 => x"39",
          2512 => x"d6",
          2513 => x"05",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"d6",
          2517 => x"05",
          2518 => x"73",
          2519 => x"38",
          2520 => x"08",
          2521 => x"53",
          2522 => x"27",
          2523 => x"d6",
          2524 => x"05",
          2525 => x"51",
          2526 => x"d6",
          2527 => x"05",
          2528 => x"e4",
          2529 => x"33",
          2530 => x"53",
          2531 => x"e4",
          2532 => x"34",
          2533 => x"08",
          2534 => x"53",
          2535 => x"ad",
          2536 => x"e4",
          2537 => x"33",
          2538 => x"53",
          2539 => x"e4",
          2540 => x"34",
          2541 => x"08",
          2542 => x"53",
          2543 => x"8d",
          2544 => x"82",
          2545 => x"ec",
          2546 => x"98",
          2547 => x"e4",
          2548 => x"33",
          2549 => x"08",
          2550 => x"54",
          2551 => x"26",
          2552 => x"0b",
          2553 => x"08",
          2554 => x"80",
          2555 => x"d6",
          2556 => x"05",
          2557 => x"d6",
          2558 => x"05",
          2559 => x"d6",
          2560 => x"05",
          2561 => x"82",
          2562 => x"fc",
          2563 => x"d6",
          2564 => x"05",
          2565 => x"81",
          2566 => x"70",
          2567 => x"52",
          2568 => x"33",
          2569 => x"08",
          2570 => x"fe",
          2571 => x"d6",
          2572 => x"05",
          2573 => x"80",
          2574 => x"82",
          2575 => x"fc",
          2576 => x"82",
          2577 => x"fc",
          2578 => x"d6",
          2579 => x"05",
          2580 => x"e4",
          2581 => x"08",
          2582 => x"81",
          2583 => x"e4",
          2584 => x"0c",
          2585 => x"08",
          2586 => x"82",
          2587 => x"8b",
          2588 => x"d6",
          2589 => x"82",
          2590 => x"02",
          2591 => x"0c",
          2592 => x"80",
          2593 => x"e4",
          2594 => x"34",
          2595 => x"08",
          2596 => x"53",
          2597 => x"82",
          2598 => x"88",
          2599 => x"08",
          2600 => x"33",
          2601 => x"d6",
          2602 => x"05",
          2603 => x"ff",
          2604 => x"a0",
          2605 => x"06",
          2606 => x"d6",
          2607 => x"05",
          2608 => x"81",
          2609 => x"53",
          2610 => x"d6",
          2611 => x"05",
          2612 => x"ad",
          2613 => x"06",
          2614 => x"0b",
          2615 => x"08",
          2616 => x"82",
          2617 => x"88",
          2618 => x"08",
          2619 => x"0c",
          2620 => x"53",
          2621 => x"d6",
          2622 => x"05",
          2623 => x"e4",
          2624 => x"33",
          2625 => x"2e",
          2626 => x"81",
          2627 => x"d6",
          2628 => x"05",
          2629 => x"81",
          2630 => x"70",
          2631 => x"72",
          2632 => x"e4",
          2633 => x"34",
          2634 => x"08",
          2635 => x"82",
          2636 => x"e8",
          2637 => x"d6",
          2638 => x"05",
          2639 => x"2e",
          2640 => x"d6",
          2641 => x"05",
          2642 => x"2e",
          2643 => x"cd",
          2644 => x"82",
          2645 => x"f4",
          2646 => x"d6",
          2647 => x"05",
          2648 => x"81",
          2649 => x"70",
          2650 => x"72",
          2651 => x"e4",
          2652 => x"34",
          2653 => x"82",
          2654 => x"e4",
          2655 => x"34",
          2656 => x"08",
          2657 => x"70",
          2658 => x"71",
          2659 => x"51",
          2660 => x"82",
          2661 => x"f8",
          2662 => x"fe",
          2663 => x"e4",
          2664 => x"33",
          2665 => x"26",
          2666 => x"0b",
          2667 => x"08",
          2668 => x"83",
          2669 => x"d6",
          2670 => x"05",
          2671 => x"73",
          2672 => x"82",
          2673 => x"f8",
          2674 => x"72",
          2675 => x"38",
          2676 => x"0b",
          2677 => x"08",
          2678 => x"82",
          2679 => x"0b",
          2680 => x"08",
          2681 => x"b2",
          2682 => x"e4",
          2683 => x"33",
          2684 => x"27",
          2685 => x"d6",
          2686 => x"05",
          2687 => x"b9",
          2688 => x"8d",
          2689 => x"82",
          2690 => x"ec",
          2691 => x"a5",
          2692 => x"82",
          2693 => x"f4",
          2694 => x"0b",
          2695 => x"08",
          2696 => x"82",
          2697 => x"f8",
          2698 => x"a0",
          2699 => x"cf",
          2700 => x"e4",
          2701 => x"33",
          2702 => x"73",
          2703 => x"82",
          2704 => x"f8",
          2705 => x"11",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"d6",
          2709 => x"05",
          2710 => x"51",
          2711 => x"d6",
          2712 => x"05",
          2713 => x"e4",
          2714 => x"33",
          2715 => x"27",
          2716 => x"d6",
          2717 => x"05",
          2718 => x"51",
          2719 => x"d6",
          2720 => x"05",
          2721 => x"e4",
          2722 => x"33",
          2723 => x"26",
          2724 => x"0b",
          2725 => x"08",
          2726 => x"81",
          2727 => x"d6",
          2728 => x"05",
          2729 => x"e4",
          2730 => x"33",
          2731 => x"74",
          2732 => x"80",
          2733 => x"e4",
          2734 => x"0c",
          2735 => x"82",
          2736 => x"f4",
          2737 => x"82",
          2738 => x"fc",
          2739 => x"82",
          2740 => x"f8",
          2741 => x"12",
          2742 => x"08",
          2743 => x"82",
          2744 => x"88",
          2745 => x"08",
          2746 => x"0c",
          2747 => x"51",
          2748 => x"72",
          2749 => x"e4",
          2750 => x"34",
          2751 => x"82",
          2752 => x"f0",
          2753 => x"72",
          2754 => x"38",
          2755 => x"08",
          2756 => x"30",
          2757 => x"08",
          2758 => x"82",
          2759 => x"8c",
          2760 => x"d6",
          2761 => x"05",
          2762 => x"53",
          2763 => x"d6",
          2764 => x"05",
          2765 => x"e4",
          2766 => x"08",
          2767 => x"0c",
          2768 => x"82",
          2769 => x"04",
          2770 => x"7a",
          2771 => x"56",
          2772 => x"80",
          2773 => x"38",
          2774 => x"15",
          2775 => x"16",
          2776 => x"d2",
          2777 => x"54",
          2778 => x"09",
          2779 => x"38",
          2780 => x"f1",
          2781 => x"76",
          2782 => x"d0",
          2783 => x"08",
          2784 => x"81",
          2785 => x"d8",
          2786 => x"d8",
          2787 => x"53",
          2788 => x"58",
          2789 => x"82",
          2790 => x"8b",
          2791 => x"33",
          2792 => x"2e",
          2793 => x"81",
          2794 => x"ff",
          2795 => x"99",
          2796 => x"38",
          2797 => x"82",
          2798 => x"8a",
          2799 => x"ff",
          2800 => x"52",
          2801 => x"81",
          2802 => x"84",
          2803 => x"dc",
          2804 => x"08",
          2805 => x"cc",
          2806 => x"39",
          2807 => x"51",
          2808 => x"82",
          2809 => x"80",
          2810 => x"b2",
          2811 => x"eb",
          2812 => x"88",
          2813 => x"39",
          2814 => x"51",
          2815 => x"82",
          2816 => x"80",
          2817 => x"b3",
          2818 => x"cf",
          2819 => x"d4",
          2820 => x"39",
          2821 => x"51",
          2822 => x"82",
          2823 => x"bb",
          2824 => x"a0",
          2825 => x"82",
          2826 => x"af",
          2827 => x"dc",
          2828 => x"82",
          2829 => x"a3",
          2830 => x"8c",
          2831 => x"82",
          2832 => x"97",
          2833 => x"b4",
          2834 => x"82",
          2835 => x"8b",
          2836 => x"e4",
          2837 => x"82",
          2838 => x"d7",
          2839 => x"3d",
          2840 => x"3d",
          2841 => x"56",
          2842 => x"e7",
          2843 => x"74",
          2844 => x"e8",
          2845 => x"39",
          2846 => x"74",
          2847 => x"3f",
          2848 => x"08",
          2849 => x"ef",
          2850 => x"d6",
          2851 => x"79",
          2852 => x"82",
          2853 => x"ff",
          2854 => x"87",
          2855 => x"ec",
          2856 => x"02",
          2857 => x"e3",
          2858 => x"57",
          2859 => x"30",
          2860 => x"73",
          2861 => x"59",
          2862 => x"77",
          2863 => x"83",
          2864 => x"74",
          2865 => x"81",
          2866 => x"55",
          2867 => x"81",
          2868 => x"53",
          2869 => x"3d",
          2870 => x"81",
          2871 => x"82",
          2872 => x"57",
          2873 => x"08",
          2874 => x"d6",
          2875 => x"c0",
          2876 => x"82",
          2877 => x"59",
          2878 => x"05",
          2879 => x"53",
          2880 => x"51",
          2881 => x"3f",
          2882 => x"08",
          2883 => x"d8",
          2884 => x"7a",
          2885 => x"2e",
          2886 => x"19",
          2887 => x"59",
          2888 => x"3d",
          2889 => x"81",
          2890 => x"76",
          2891 => x"07",
          2892 => x"30",
          2893 => x"72",
          2894 => x"51",
          2895 => x"2e",
          2896 => x"b6",
          2897 => x"c0",
          2898 => x"52",
          2899 => x"92",
          2900 => x"75",
          2901 => x"0c",
          2902 => x"04",
          2903 => x"7d",
          2904 => x"bb",
          2905 => x"5a",
          2906 => x"53",
          2907 => x"51",
          2908 => x"82",
          2909 => x"80",
          2910 => x"80",
          2911 => x"77",
          2912 => x"38",
          2913 => x"f2",
          2914 => x"f2",
          2915 => x"f2",
          2916 => x"f2",
          2917 => x"82",
          2918 => x"53",
          2919 => x"08",
          2920 => x"ac",
          2921 => x"b0",
          2922 => x"b8",
          2923 => x"61",
          2924 => x"d8",
          2925 => x"7f",
          2926 => x"82",
          2927 => x"59",
          2928 => x"04",
          2929 => x"d8",
          2930 => x"0d",
          2931 => x"0d",
          2932 => x"02",
          2933 => x"cf",
          2934 => x"73",
          2935 => x"5f",
          2936 => x"5e",
          2937 => x"82",
          2938 => x"ff",
          2939 => x"82",
          2940 => x"ff",
          2941 => x"80",
          2942 => x"27",
          2943 => x"7b",
          2944 => x"38",
          2945 => x"a7",
          2946 => x"39",
          2947 => x"72",
          2948 => x"38",
          2949 => x"82",
          2950 => x"ff",
          2951 => x"89",
          2952 => x"f8",
          2953 => x"b0",
          2954 => x"55",
          2955 => x"74",
          2956 => x"7a",
          2957 => x"72",
          2958 => x"b6",
          2959 => x"b7",
          2960 => x"39",
          2961 => x"51",
          2962 => x"3f",
          2963 => x"a1",
          2964 => x"53",
          2965 => x"8e",
          2966 => x"52",
          2967 => x"51",
          2968 => x"3f",
          2969 => x"b7",
          2970 => x"b6",
          2971 => x"15",
          2972 => x"bc",
          2973 => x"51",
          2974 => x"fe",
          2975 => x"b7",
          2976 => x"b6",
          2977 => x"55",
          2978 => x"80",
          2979 => x"18",
          2980 => x"53",
          2981 => x"7a",
          2982 => x"81",
          2983 => x"9f",
          2984 => x"38",
          2985 => x"73",
          2986 => x"ff",
          2987 => x"72",
          2988 => x"38",
          2989 => x"26",
          2990 => x"f2",
          2991 => x"73",
          2992 => x"82",
          2993 => x"52",
          2994 => x"e6",
          2995 => x"55",
          2996 => x"82",
          2997 => x"d2",
          2998 => x"18",
          2999 => x"58",
          3000 => x"82",
          3001 => x"98",
          3002 => x"2c",
          3003 => x"a0",
          3004 => x"06",
          3005 => x"d1",
          3006 => x"d8",
          3007 => x"70",
          3008 => x"a0",
          3009 => x"72",
          3010 => x"30",
          3011 => x"73",
          3012 => x"51",
          3013 => x"57",
          3014 => x"73",
          3015 => x"76",
          3016 => x"81",
          3017 => x"80",
          3018 => x"7c",
          3019 => x"78",
          3020 => x"38",
          3021 => x"82",
          3022 => x"8f",
          3023 => x"fc",
          3024 => x"9b",
          3025 => x"b7",
          3026 => x"b7",
          3027 => x"ff",
          3028 => x"82",
          3029 => x"51",
          3030 => x"82",
          3031 => x"82",
          3032 => x"82",
          3033 => x"52",
          3034 => x"51",
          3035 => x"3f",
          3036 => x"84",
          3037 => x"3f",
          3038 => x"04",
          3039 => x"87",
          3040 => x"08",
          3041 => x"3f",
          3042 => x"bd",
          3043 => x"d4",
          3044 => x"3f",
          3045 => x"b1",
          3046 => x"2a",
          3047 => x"51",
          3048 => x"2e",
          3049 => x"51",
          3050 => x"82",
          3051 => x"99",
          3052 => x"51",
          3053 => x"72",
          3054 => x"81",
          3055 => x"71",
          3056 => x"38",
          3057 => x"81",
          3058 => x"fc",
          3059 => x"3f",
          3060 => x"f5",
          3061 => x"2a",
          3062 => x"51",
          3063 => x"2e",
          3064 => x"51",
          3065 => x"82",
          3066 => x"98",
          3067 => x"51",
          3068 => x"72",
          3069 => x"81",
          3070 => x"71",
          3071 => x"38",
          3072 => x"c5",
          3073 => x"a0",
          3074 => x"3f",
          3075 => x"b9",
          3076 => x"2a",
          3077 => x"51",
          3078 => x"2e",
          3079 => x"51",
          3080 => x"82",
          3081 => x"98",
          3082 => x"51",
          3083 => x"72",
          3084 => x"81",
          3085 => x"71",
          3086 => x"38",
          3087 => x"89",
          3088 => x"c8",
          3089 => x"3f",
          3090 => x"fd",
          3091 => x"2a",
          3092 => x"51",
          3093 => x"2e",
          3094 => x"51",
          3095 => x"82",
          3096 => x"97",
          3097 => x"51",
          3098 => x"72",
          3099 => x"81",
          3100 => x"71",
          3101 => x"38",
          3102 => x"cd",
          3103 => x"f0",
          3104 => x"3f",
          3105 => x"c1",
          3106 => x"3f",
          3107 => x"04",
          3108 => x"77",
          3109 => x"a3",
          3110 => x"55",
          3111 => x"52",
          3112 => x"ed",
          3113 => x"82",
          3114 => x"54",
          3115 => x"81",
          3116 => x"ac",
          3117 => x"e8",
          3118 => x"f1",
          3119 => x"d8",
          3120 => x"82",
          3121 => x"07",
          3122 => x"71",
          3123 => x"54",
          3124 => x"82",
          3125 => x"0b",
          3126 => x"c8",
          3127 => x"81",
          3128 => x"06",
          3129 => x"ed",
          3130 => x"52",
          3131 => x"c5",
          3132 => x"d6",
          3133 => x"2e",
          3134 => x"d6",
          3135 => x"cd",
          3136 => x"39",
          3137 => x"51",
          3138 => x"3f",
          3139 => x"0b",
          3140 => x"34",
          3141 => x"d0",
          3142 => x"73",
          3143 => x"81",
          3144 => x"82",
          3145 => x"74",
          3146 => x"a9",
          3147 => x"0b",
          3148 => x"0c",
          3149 => x"04",
          3150 => x"80",
          3151 => x"ff",
          3152 => x"e4",
          3153 => x"52",
          3154 => x"c8",
          3155 => x"d6",
          3156 => x"ff",
          3157 => x"7e",
          3158 => x"06",
          3159 => x"3d",
          3160 => x"82",
          3161 => x"78",
          3162 => x"3f",
          3163 => x"52",
          3164 => x"51",
          3165 => x"3f",
          3166 => x"08",
          3167 => x"38",
          3168 => x"51",
          3169 => x"81",
          3170 => x"82",
          3171 => x"ff",
          3172 => x"97",
          3173 => x"5a",
          3174 => x"79",
          3175 => x"3f",
          3176 => x"84",
          3177 => x"a0",
          3178 => x"d8",
          3179 => x"70",
          3180 => x"59",
          3181 => x"2e",
          3182 => x"78",
          3183 => x"b2",
          3184 => x"2e",
          3185 => x"78",
          3186 => x"38",
          3187 => x"ff",
          3188 => x"bc",
          3189 => x"38",
          3190 => x"78",
          3191 => x"83",
          3192 => x"80",
          3193 => x"cd",
          3194 => x"2e",
          3195 => x"8a",
          3196 => x"80",
          3197 => x"db",
          3198 => x"f9",
          3199 => x"78",
          3200 => x"88",
          3201 => x"80",
          3202 => x"a3",
          3203 => x"39",
          3204 => x"2e",
          3205 => x"78",
          3206 => x"8b",
          3207 => x"82",
          3208 => x"38",
          3209 => x"78",
          3210 => x"89",
          3211 => x"80",
          3212 => x"ff",
          3213 => x"ff",
          3214 => x"ec",
          3215 => x"d6",
          3216 => x"2e",
          3217 => x"b5",
          3218 => x"11",
          3219 => x"05",
          3220 => x"3f",
          3221 => x"08",
          3222 => x"af",
          3223 => x"fe",
          3224 => x"ff",
          3225 => x"ec",
          3226 => x"d6",
          3227 => x"38",
          3228 => x"08",
          3229 => x"84",
          3230 => x"dc",
          3231 => x"5c",
          3232 => x"27",
          3233 => x"62",
          3234 => x"70",
          3235 => x"0c",
          3236 => x"f5",
          3237 => x"39",
          3238 => x"80",
          3239 => x"84",
          3240 => x"d3",
          3241 => x"d8",
          3242 => x"fd",
          3243 => x"3d",
          3244 => x"53",
          3245 => x"51",
          3246 => x"82",
          3247 => x"80",
          3248 => x"38",
          3249 => x"f8",
          3250 => x"84",
          3251 => x"a7",
          3252 => x"d8",
          3253 => x"fd",
          3254 => x"ba",
          3255 => x"ad",
          3256 => x"5a",
          3257 => x"81",
          3258 => x"59",
          3259 => x"05",
          3260 => x"34",
          3261 => x"43",
          3262 => x"3d",
          3263 => x"53",
          3264 => x"51",
          3265 => x"82",
          3266 => x"80",
          3267 => x"38",
          3268 => x"fc",
          3269 => x"84",
          3270 => x"db",
          3271 => x"d8",
          3272 => x"fc",
          3273 => x"3d",
          3274 => x"53",
          3275 => x"51",
          3276 => x"82",
          3277 => x"80",
          3278 => x"38",
          3279 => x"51",
          3280 => x"3f",
          3281 => x"64",
          3282 => x"62",
          3283 => x"33",
          3284 => x"78",
          3285 => x"38",
          3286 => x"54",
          3287 => x"79",
          3288 => x"b0",
          3289 => x"f0",
          3290 => x"63",
          3291 => x"5a",
          3292 => x"51",
          3293 => x"fc",
          3294 => x"3d",
          3295 => x"53",
          3296 => x"51",
          3297 => x"82",
          3298 => x"80",
          3299 => x"d4",
          3300 => x"78",
          3301 => x"38",
          3302 => x"08",
          3303 => x"39",
          3304 => x"33",
          3305 => x"2e",
          3306 => x"d3",
          3307 => x"bc",
          3308 => x"ba",
          3309 => x"80",
          3310 => x"82",
          3311 => x"45",
          3312 => x"d4",
          3313 => x"78",
          3314 => x"38",
          3315 => x"08",
          3316 => x"82",
          3317 => x"59",
          3318 => x"88",
          3319 => x"90",
          3320 => x"39",
          3321 => x"08",
          3322 => x"45",
          3323 => x"fc",
          3324 => x"84",
          3325 => x"ff",
          3326 => x"d8",
          3327 => x"38",
          3328 => x"33",
          3329 => x"2e",
          3330 => x"d3",
          3331 => x"80",
          3332 => x"d4",
          3333 => x"78",
          3334 => x"38",
          3335 => x"08",
          3336 => x"82",
          3337 => x"59",
          3338 => x"88",
          3339 => x"84",
          3340 => x"39",
          3341 => x"33",
          3342 => x"2e",
          3343 => x"d4",
          3344 => x"99",
          3345 => x"b6",
          3346 => x"80",
          3347 => x"82",
          3348 => x"44",
          3349 => x"d4",
          3350 => x"05",
          3351 => x"fe",
          3352 => x"ff",
          3353 => x"e8",
          3354 => x"d6",
          3355 => x"2e",
          3356 => x"63",
          3357 => x"88",
          3358 => x"81",
          3359 => x"32",
          3360 => x"72",
          3361 => x"70",
          3362 => x"51",
          3363 => x"80",
          3364 => x"7a",
          3365 => x"38",
          3366 => x"ba",
          3367 => x"c3",
          3368 => x"64",
          3369 => x"63",
          3370 => x"f2",
          3371 => x"ba",
          3372 => x"b1",
          3373 => x"ff",
          3374 => x"ff",
          3375 => x"e7",
          3376 => x"d6",
          3377 => x"2e",
          3378 => x"b5",
          3379 => x"11",
          3380 => x"05",
          3381 => x"3f",
          3382 => x"08",
          3383 => x"38",
          3384 => x"80",
          3385 => x"79",
          3386 => x"05",
          3387 => x"fe",
          3388 => x"ff",
          3389 => x"e6",
          3390 => x"d6",
          3391 => x"38",
          3392 => x"64",
          3393 => x"52",
          3394 => x"51",
          3395 => x"3f",
          3396 => x"08",
          3397 => x"52",
          3398 => x"aa",
          3399 => x"46",
          3400 => x"78",
          3401 => x"e3",
          3402 => x"27",
          3403 => x"3d",
          3404 => x"53",
          3405 => x"51",
          3406 => x"82",
          3407 => x"80",
          3408 => x"64",
          3409 => x"cf",
          3410 => x"34",
          3411 => x"45",
          3412 => x"82",
          3413 => x"c5",
          3414 => x"a7",
          3415 => x"fe",
          3416 => x"ff",
          3417 => x"e0",
          3418 => x"d6",
          3419 => x"2e",
          3420 => x"b5",
          3421 => x"11",
          3422 => x"05",
          3423 => x"3f",
          3424 => x"08",
          3425 => x"38",
          3426 => x"80",
          3427 => x"79",
          3428 => x"5b",
          3429 => x"b5",
          3430 => x"11",
          3431 => x"05",
          3432 => x"3f",
          3433 => x"08",
          3434 => x"df",
          3435 => x"22",
          3436 => x"ba",
          3437 => x"a8",
          3438 => x"f2",
          3439 => x"80",
          3440 => x"51",
          3441 => x"3f",
          3442 => x"33",
          3443 => x"2e",
          3444 => x"78",
          3445 => x"38",
          3446 => x"42",
          3447 => x"3d",
          3448 => x"53",
          3449 => x"51",
          3450 => x"82",
          3451 => x"80",
          3452 => x"61",
          3453 => x"c2",
          3454 => x"70",
          3455 => x"23",
          3456 => x"a9",
          3457 => x"f0",
          3458 => x"3f",
          3459 => x"b5",
          3460 => x"11",
          3461 => x"05",
          3462 => x"3f",
          3463 => x"08",
          3464 => x"e7",
          3465 => x"fe",
          3466 => x"ff",
          3467 => x"de",
          3468 => x"d6",
          3469 => x"2e",
          3470 => x"61",
          3471 => x"61",
          3472 => x"b5",
          3473 => x"11",
          3474 => x"05",
          3475 => x"3f",
          3476 => x"08",
          3477 => x"b3",
          3478 => x"08",
          3479 => x"bb",
          3480 => x"a6",
          3481 => x"f2",
          3482 => x"80",
          3483 => x"51",
          3484 => x"3f",
          3485 => x"33",
          3486 => x"2e",
          3487 => x"9f",
          3488 => x"38",
          3489 => x"f0",
          3490 => x"84",
          3491 => x"96",
          3492 => x"d8",
          3493 => x"8d",
          3494 => x"71",
          3495 => x"84",
          3496 => x"b5",
          3497 => x"f0",
          3498 => x"3f",
          3499 => x"b5",
          3500 => x"11",
          3501 => x"05",
          3502 => x"3f",
          3503 => x"08",
          3504 => x"c7",
          3505 => x"82",
          3506 => x"ff",
          3507 => x"64",
          3508 => x"b5",
          3509 => x"11",
          3510 => x"05",
          3511 => x"3f",
          3512 => x"08",
          3513 => x"a3",
          3514 => x"82",
          3515 => x"ff",
          3516 => x"64",
          3517 => x"82",
          3518 => x"80",
          3519 => x"38",
          3520 => x"08",
          3521 => x"c8",
          3522 => x"cc",
          3523 => x"39",
          3524 => x"51",
          3525 => x"ff",
          3526 => x"f4",
          3527 => x"bc",
          3528 => x"bf",
          3529 => x"ff",
          3530 => x"bf",
          3531 => x"39",
          3532 => x"59",
          3533 => x"f4",
          3534 => x"f8",
          3535 => x"d2",
          3536 => x"d6",
          3537 => x"82",
          3538 => x"80",
          3539 => x"38",
          3540 => x"08",
          3541 => x"ff",
          3542 => x"84",
          3543 => x"d6",
          3544 => x"7f",
          3545 => x"78",
          3546 => x"d2",
          3547 => x"d8",
          3548 => x"91",
          3549 => x"d8",
          3550 => x"81",
          3551 => x"5b",
          3552 => x"b2",
          3553 => x"24",
          3554 => x"81",
          3555 => x"80",
          3556 => x"83",
          3557 => x"80",
          3558 => x"bc",
          3559 => x"55",
          3560 => x"54",
          3561 => x"bc",
          3562 => x"3d",
          3563 => x"51",
          3564 => x"3f",
          3565 => x"52",
          3566 => x"b0",
          3567 => x"b3",
          3568 => x"7b",
          3569 => x"98",
          3570 => x"82",
          3571 => x"b5",
          3572 => x"05",
          3573 => x"e8",
          3574 => x"7b",
          3575 => x"82",
          3576 => x"b5",
          3577 => x"05",
          3578 => x"d4",
          3579 => x"f0",
          3580 => x"88",
          3581 => x"65",
          3582 => x"84",
          3583 => x"84",
          3584 => x"b5",
          3585 => x"05",
          3586 => x"3f",
          3587 => x"08",
          3588 => x"08",
          3589 => x"70",
          3590 => x"25",
          3591 => x"5f",
          3592 => x"83",
          3593 => x"81",
          3594 => x"06",
          3595 => x"2e",
          3596 => x"1b",
          3597 => x"06",
          3598 => x"fe",
          3599 => x"81",
          3600 => x"32",
          3601 => x"89",
          3602 => x"2e",
          3603 => x"89",
          3604 => x"c0",
          3605 => x"8b",
          3606 => x"b1",
          3607 => x"ab",
          3608 => x"d0",
          3609 => x"fb",
          3610 => x"39",
          3611 => x"80",
          3612 => x"88",
          3613 => x"94",
          3614 => x"87",
          3615 => x"72",
          3616 => x"3f",
          3617 => x"08",
          3618 => x"c0",
          3619 => x"55",
          3620 => x"80",
          3621 => x"d7",
          3622 => x"82",
          3623 => x"07",
          3624 => x"8c",
          3625 => x"94",
          3626 => x"87",
          3627 => x"72",
          3628 => x"3f",
          3629 => x"08",
          3630 => x"c0",
          3631 => x"55",
          3632 => x"80",
          3633 => x"d6",
          3634 => x"82",
          3635 => x"07",
          3636 => x"9c",
          3637 => x"83",
          3638 => x"94",
          3639 => x"80",
          3640 => x"c0",
          3641 => x"87",
          3642 => x"53",
          3643 => x"84",
          3644 => x"87",
          3645 => x"73",
          3646 => x"87",
          3647 => x"53",
          3648 => x"e2",
          3649 => x"84",
          3650 => x"87",
          3651 => x"73",
          3652 => x"80",
          3653 => x"51",
          3654 => x"80",
          3655 => x"51",
          3656 => x"80",
          3657 => x"51",
          3658 => x"80",
          3659 => x"51",
          3660 => x"80",
          3661 => x"51",
          3662 => x"80",
          3663 => x"a6",
          3664 => x"52",
          3665 => x"f0",
          3666 => x"b8",
          3667 => x"ca",
          3668 => x"84",
          3669 => x"34",
          3670 => x"3d",
          3671 => x"c0",
          3672 => x"f2",
          3673 => x"f2",
          3674 => x"bc",
          3675 => x"bc",
          3676 => x"ab",
          3677 => x"3f",
          3678 => x"51",
          3679 => x"3f",
          3680 => x"51",
          3681 => x"3f",
          3682 => x"51",
          3683 => x"81",
          3684 => x"3f",
          3685 => x"80",
          3686 => x"0d",
          3687 => x"53",
          3688 => x"52",
          3689 => x"82",
          3690 => x"81",
          3691 => x"07",
          3692 => x"52",
          3693 => x"e8",
          3694 => x"d6",
          3695 => x"3d",
          3696 => x"3d",
          3697 => x"08",
          3698 => x"73",
          3699 => x"74",
          3700 => x"38",
          3701 => x"70",
          3702 => x"81",
          3703 => x"81",
          3704 => x"39",
          3705 => x"70",
          3706 => x"81",
          3707 => x"81",
          3708 => x"54",
          3709 => x"81",
          3710 => x"06",
          3711 => x"39",
          3712 => x"80",
          3713 => x"54",
          3714 => x"83",
          3715 => x"70",
          3716 => x"38",
          3717 => x"98",
          3718 => x"52",
          3719 => x"52",
          3720 => x"2e",
          3721 => x"54",
          3722 => x"84",
          3723 => x"38",
          3724 => x"52",
          3725 => x"2e",
          3726 => x"83",
          3727 => x"70",
          3728 => x"30",
          3729 => x"76",
          3730 => x"51",
          3731 => x"88",
          3732 => x"70",
          3733 => x"34",
          3734 => x"72",
          3735 => x"d6",
          3736 => x"3d",
          3737 => x"3d",
          3738 => x"72",
          3739 => x"91",
          3740 => x"fc",
          3741 => x"51",
          3742 => x"82",
          3743 => x"85",
          3744 => x"83",
          3745 => x"72",
          3746 => x"0c",
          3747 => x"04",
          3748 => x"76",
          3749 => x"ff",
          3750 => x"81",
          3751 => x"26",
          3752 => x"83",
          3753 => x"05",
          3754 => x"70",
          3755 => x"8a",
          3756 => x"33",
          3757 => x"70",
          3758 => x"fe",
          3759 => x"33",
          3760 => x"70",
          3761 => x"f2",
          3762 => x"33",
          3763 => x"70",
          3764 => x"e6",
          3765 => x"22",
          3766 => x"74",
          3767 => x"80",
          3768 => x"13",
          3769 => x"52",
          3770 => x"26",
          3771 => x"81",
          3772 => x"98",
          3773 => x"22",
          3774 => x"bc",
          3775 => x"33",
          3776 => x"b8",
          3777 => x"33",
          3778 => x"b4",
          3779 => x"33",
          3780 => x"b0",
          3781 => x"33",
          3782 => x"ac",
          3783 => x"33",
          3784 => x"a8",
          3785 => x"c0",
          3786 => x"73",
          3787 => x"a0",
          3788 => x"87",
          3789 => x"0c",
          3790 => x"82",
          3791 => x"86",
          3792 => x"f3",
          3793 => x"5b",
          3794 => x"9c",
          3795 => x"0c",
          3796 => x"bc",
          3797 => x"7b",
          3798 => x"98",
          3799 => x"79",
          3800 => x"87",
          3801 => x"08",
          3802 => x"1c",
          3803 => x"98",
          3804 => x"79",
          3805 => x"87",
          3806 => x"08",
          3807 => x"1c",
          3808 => x"98",
          3809 => x"79",
          3810 => x"87",
          3811 => x"08",
          3812 => x"1c",
          3813 => x"98",
          3814 => x"79",
          3815 => x"80",
          3816 => x"83",
          3817 => x"59",
          3818 => x"ff",
          3819 => x"1b",
          3820 => x"1b",
          3821 => x"1b",
          3822 => x"1b",
          3823 => x"1b",
          3824 => x"83",
          3825 => x"52",
          3826 => x"51",
          3827 => x"3f",
          3828 => x"04",
          3829 => x"02",
          3830 => x"82",
          3831 => x"70",
          3832 => x"58",
          3833 => x"c0",
          3834 => x"75",
          3835 => x"38",
          3836 => x"94",
          3837 => x"70",
          3838 => x"81",
          3839 => x"52",
          3840 => x"8c",
          3841 => x"2a",
          3842 => x"51",
          3843 => x"38",
          3844 => x"70",
          3845 => x"51",
          3846 => x"8d",
          3847 => x"2a",
          3848 => x"51",
          3849 => x"be",
          3850 => x"ff",
          3851 => x"c0",
          3852 => x"70",
          3853 => x"38",
          3854 => x"90",
          3855 => x"0c",
          3856 => x"d8",
          3857 => x"0d",
          3858 => x"0d",
          3859 => x"33",
          3860 => x"9f",
          3861 => x"52",
          3862 => x"ec",
          3863 => x"0d",
          3864 => x"0d",
          3865 => x"74",
          3866 => x"ff",
          3867 => x"57",
          3868 => x"80",
          3869 => x"81",
          3870 => x"15",
          3871 => x"33",
          3872 => x"06",
          3873 => x"58",
          3874 => x"84",
          3875 => x"2e",
          3876 => x"c0",
          3877 => x"70",
          3878 => x"2a",
          3879 => x"53",
          3880 => x"80",
          3881 => x"71",
          3882 => x"81",
          3883 => x"70",
          3884 => x"81",
          3885 => x"06",
          3886 => x"80",
          3887 => x"71",
          3888 => x"81",
          3889 => x"70",
          3890 => x"74",
          3891 => x"51",
          3892 => x"80",
          3893 => x"2e",
          3894 => x"c0",
          3895 => x"77",
          3896 => x"17",
          3897 => x"81",
          3898 => x"53",
          3899 => x"86",
          3900 => x"d6",
          3901 => x"3d",
          3902 => x"3d",
          3903 => x"ec",
          3904 => x"ff",
          3905 => x"87",
          3906 => x"51",
          3907 => x"86",
          3908 => x"94",
          3909 => x"08",
          3910 => x"70",
          3911 => x"51",
          3912 => x"2e",
          3913 => x"81",
          3914 => x"87",
          3915 => x"52",
          3916 => x"86",
          3917 => x"94",
          3918 => x"08",
          3919 => x"06",
          3920 => x"0c",
          3921 => x"0d",
          3922 => x"0d",
          3923 => x"33",
          3924 => x"06",
          3925 => x"c0",
          3926 => x"70",
          3927 => x"38",
          3928 => x"94",
          3929 => x"70",
          3930 => x"81",
          3931 => x"51",
          3932 => x"80",
          3933 => x"72",
          3934 => x"51",
          3935 => x"80",
          3936 => x"2e",
          3937 => x"c0",
          3938 => x"71",
          3939 => x"2b",
          3940 => x"51",
          3941 => x"82",
          3942 => x"84",
          3943 => x"ff",
          3944 => x"c0",
          3945 => x"70",
          3946 => x"06",
          3947 => x"80",
          3948 => x"38",
          3949 => x"a4",
          3950 => x"f0",
          3951 => x"9e",
          3952 => x"d3",
          3953 => x"c0",
          3954 => x"82",
          3955 => x"87",
          3956 => x"08",
          3957 => x"0c",
          3958 => x"9c",
          3959 => x"80",
          3960 => x"9e",
          3961 => x"d4",
          3962 => x"c0",
          3963 => x"82",
          3964 => x"87",
          3965 => x"08",
          3966 => x"0c",
          3967 => x"b4",
          3968 => x"90",
          3969 => x"9e",
          3970 => x"d4",
          3971 => x"c0",
          3972 => x"82",
          3973 => x"87",
          3974 => x"08",
          3975 => x"0c",
          3976 => x"c4",
          3977 => x"a0",
          3978 => x"9e",
          3979 => x"70",
          3980 => x"23",
          3981 => x"84",
          3982 => x"a8",
          3983 => x"9e",
          3984 => x"d4",
          3985 => x"c0",
          3986 => x"82",
          3987 => x"81",
          3988 => x"b4",
          3989 => x"87",
          3990 => x"08",
          3991 => x"0a",
          3992 => x"52",
          3993 => x"83",
          3994 => x"71",
          3995 => x"34",
          3996 => x"c0",
          3997 => x"70",
          3998 => x"06",
          3999 => x"70",
          4000 => x"38",
          4001 => x"82",
          4002 => x"80",
          4003 => x"9e",
          4004 => x"90",
          4005 => x"51",
          4006 => x"80",
          4007 => x"81",
          4008 => x"d4",
          4009 => x"0b",
          4010 => x"90",
          4011 => x"80",
          4012 => x"52",
          4013 => x"2e",
          4014 => x"52",
          4015 => x"b8",
          4016 => x"87",
          4017 => x"08",
          4018 => x"80",
          4019 => x"52",
          4020 => x"83",
          4021 => x"71",
          4022 => x"34",
          4023 => x"c0",
          4024 => x"70",
          4025 => x"06",
          4026 => x"70",
          4027 => x"38",
          4028 => x"82",
          4029 => x"80",
          4030 => x"9e",
          4031 => x"84",
          4032 => x"51",
          4033 => x"80",
          4034 => x"81",
          4035 => x"d4",
          4036 => x"0b",
          4037 => x"90",
          4038 => x"80",
          4039 => x"52",
          4040 => x"2e",
          4041 => x"52",
          4042 => x"bc",
          4043 => x"87",
          4044 => x"08",
          4045 => x"80",
          4046 => x"52",
          4047 => x"83",
          4048 => x"71",
          4049 => x"34",
          4050 => x"c0",
          4051 => x"70",
          4052 => x"06",
          4053 => x"70",
          4054 => x"38",
          4055 => x"82",
          4056 => x"80",
          4057 => x"9e",
          4058 => x"a0",
          4059 => x"52",
          4060 => x"2e",
          4061 => x"52",
          4062 => x"bf",
          4063 => x"9e",
          4064 => x"98",
          4065 => x"8a",
          4066 => x"51",
          4067 => x"c0",
          4068 => x"87",
          4069 => x"08",
          4070 => x"06",
          4071 => x"70",
          4072 => x"38",
          4073 => x"82",
          4074 => x"87",
          4075 => x"08",
          4076 => x"06",
          4077 => x"51",
          4078 => x"82",
          4079 => x"80",
          4080 => x"9e",
          4081 => x"88",
          4082 => x"52",
          4083 => x"83",
          4084 => x"71",
          4085 => x"34",
          4086 => x"90",
          4087 => x"06",
          4088 => x"82",
          4089 => x"83",
          4090 => x"fb",
          4091 => x"bd",
          4092 => x"93",
          4093 => x"d4",
          4094 => x"73",
          4095 => x"38",
          4096 => x"51",
          4097 => x"3f",
          4098 => x"51",
          4099 => x"3f",
          4100 => x"33",
          4101 => x"2e",
          4102 => x"d4",
          4103 => x"d4",
          4104 => x"54",
          4105 => x"88",
          4106 => x"ac",
          4107 => x"bb",
          4108 => x"80",
          4109 => x"82",
          4110 => x"82",
          4111 => x"11",
          4112 => x"be",
          4113 => x"93",
          4114 => x"d4",
          4115 => x"73",
          4116 => x"38",
          4117 => x"08",
          4118 => x"08",
          4119 => x"82",
          4120 => x"ff",
          4121 => x"82",
          4122 => x"54",
          4123 => x"94",
          4124 => x"f8",
          4125 => x"fc",
          4126 => x"52",
          4127 => x"51",
          4128 => x"3f",
          4129 => x"33",
          4130 => x"2e",
          4131 => x"d4",
          4132 => x"d4",
          4133 => x"54",
          4134 => x"f8",
          4135 => x"b8",
          4136 => x"bf",
          4137 => x"80",
          4138 => x"82",
          4139 => x"52",
          4140 => x"51",
          4141 => x"3f",
          4142 => x"33",
          4143 => x"2e",
          4144 => x"d4",
          4145 => x"82",
          4146 => x"ff",
          4147 => x"82",
          4148 => x"54",
          4149 => x"8e",
          4150 => x"c2",
          4151 => x"bf",
          4152 => x"91",
          4153 => x"d4",
          4154 => x"73",
          4155 => x"38",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"33",
          4159 => x"2e",
          4160 => x"c0",
          4161 => x"ad",
          4162 => x"d4",
          4163 => x"73",
          4164 => x"38",
          4165 => x"51",
          4166 => x"3f",
          4167 => x"33",
          4168 => x"2e",
          4169 => x"c0",
          4170 => x"ad",
          4171 => x"d4",
          4172 => x"73",
          4173 => x"38",
          4174 => x"51",
          4175 => x"3f",
          4176 => x"51",
          4177 => x"3f",
          4178 => x"08",
          4179 => x"bc",
          4180 => x"84",
          4181 => x"9c",
          4182 => x"c0",
          4183 => x"90",
          4184 => x"d4",
          4185 => x"82",
          4186 => x"ff",
          4187 => x"82",
          4188 => x"ff",
          4189 => x"82",
          4190 => x"52",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"08",
          4194 => x"c0",
          4195 => x"c5",
          4196 => x"d6",
          4197 => x"84",
          4198 => x"71",
          4199 => x"82",
          4200 => x"52",
          4201 => x"51",
          4202 => x"3f",
          4203 => x"33",
          4204 => x"2e",
          4205 => x"d4",
          4206 => x"bd",
          4207 => x"75",
          4208 => x"3f",
          4209 => x"08",
          4210 => x"29",
          4211 => x"54",
          4212 => x"d8",
          4213 => x"c2",
          4214 => x"8f",
          4215 => x"d4",
          4216 => x"73",
          4217 => x"38",
          4218 => x"08",
          4219 => x"c0",
          4220 => x"c4",
          4221 => x"d6",
          4222 => x"84",
          4223 => x"71",
          4224 => x"82",
          4225 => x"52",
          4226 => x"51",
          4227 => x"3f",
          4228 => x"ae",
          4229 => x"3d",
          4230 => x"3d",
          4231 => x"05",
          4232 => x"52",
          4233 => x"aa",
          4234 => x"29",
          4235 => x"05",
          4236 => x"04",
          4237 => x"51",
          4238 => x"c2",
          4239 => x"39",
          4240 => x"51",
          4241 => x"c3",
          4242 => x"39",
          4243 => x"51",
          4244 => x"c3",
          4245 => x"8e",
          4246 => x"3d",
          4247 => x"88",
          4248 => x"80",
          4249 => x"96",
          4250 => x"82",
          4251 => x"87",
          4252 => x"0c",
          4253 => x"0d",
          4254 => x"70",
          4255 => x"98",
          4256 => x"2c",
          4257 => x"70",
          4258 => x"53",
          4259 => x"51",
          4260 => x"c3",
          4261 => x"55",
          4262 => x"25",
          4263 => x"c3",
          4264 => x"12",
          4265 => x"97",
          4266 => x"33",
          4267 => x"70",
          4268 => x"81",
          4269 => x"81",
          4270 => x"d6",
          4271 => x"3d",
          4272 => x"3d",
          4273 => x"84",
          4274 => x"33",
          4275 => x"56",
          4276 => x"2e",
          4277 => x"f2",
          4278 => x"88",
          4279 => x"d2",
          4280 => x"bc",
          4281 => x"51",
          4282 => x"3f",
          4283 => x"08",
          4284 => x"ff",
          4285 => x"73",
          4286 => x"53",
          4287 => x"72",
          4288 => x"53",
          4289 => x"51",
          4290 => x"3f",
          4291 => x"87",
          4292 => x"f6",
          4293 => x"02",
          4294 => x"05",
          4295 => x"05",
          4296 => x"82",
          4297 => x"70",
          4298 => x"d4",
          4299 => x"08",
          4300 => x"5a",
          4301 => x"80",
          4302 => x"74",
          4303 => x"3f",
          4304 => x"33",
          4305 => x"82",
          4306 => x"81",
          4307 => x"58",
          4308 => x"94",
          4309 => x"d8",
          4310 => x"82",
          4311 => x"70",
          4312 => x"d4",
          4313 => x"08",
          4314 => x"74",
          4315 => x"38",
          4316 => x"52",
          4317 => x"b6",
          4318 => x"d5",
          4319 => x"05",
          4320 => x"d5",
          4321 => x"81",
          4322 => x"93",
          4323 => x"38",
          4324 => x"d5",
          4325 => x"80",
          4326 => x"82",
          4327 => x"56",
          4328 => x"ac",
          4329 => x"9c",
          4330 => x"a4",
          4331 => x"fc",
          4332 => x"53",
          4333 => x"51",
          4334 => x"3f",
          4335 => x"08",
          4336 => x"81",
          4337 => x"82",
          4338 => x"51",
          4339 => x"3f",
          4340 => x"04",
          4341 => x"82",
          4342 => x"93",
          4343 => x"52",
          4344 => x"89",
          4345 => x"9a",
          4346 => x"73",
          4347 => x"84",
          4348 => x"73",
          4349 => x"38",
          4350 => x"d5",
          4351 => x"d5",
          4352 => x"71",
          4353 => x"38",
          4354 => x"f1",
          4355 => x"d5",
          4356 => x"9a",
          4357 => x"0b",
          4358 => x"0c",
          4359 => x"04",
          4360 => x"81",
          4361 => x"82",
          4362 => x"51",
          4363 => x"3f",
          4364 => x"08",
          4365 => x"82",
          4366 => x"53",
          4367 => x"88",
          4368 => x"56",
          4369 => x"3f",
          4370 => x"08",
          4371 => x"38",
          4372 => x"b3",
          4373 => x"d6",
          4374 => x"80",
          4375 => x"d8",
          4376 => x"38",
          4377 => x"08",
          4378 => x"17",
          4379 => x"74",
          4380 => x"76",
          4381 => x"82",
          4382 => x"57",
          4383 => x"3f",
          4384 => x"09",
          4385 => x"af",
          4386 => x"0d",
          4387 => x"0d",
          4388 => x"ad",
          4389 => x"5a",
          4390 => x"58",
          4391 => x"d5",
          4392 => x"80",
          4393 => x"82",
          4394 => x"81",
          4395 => x"0b",
          4396 => x"08",
          4397 => x"f8",
          4398 => x"70",
          4399 => x"9d",
          4400 => x"d6",
          4401 => x"2e",
          4402 => x"51",
          4403 => x"3f",
          4404 => x"08",
          4405 => x"55",
          4406 => x"d6",
          4407 => x"8e",
          4408 => x"d8",
          4409 => x"70",
          4410 => x"80",
          4411 => x"09",
          4412 => x"72",
          4413 => x"51",
          4414 => x"77",
          4415 => x"73",
          4416 => x"82",
          4417 => x"8c",
          4418 => x"51",
          4419 => x"3f",
          4420 => x"08",
          4421 => x"38",
          4422 => x"51",
          4423 => x"3f",
          4424 => x"09",
          4425 => x"38",
          4426 => x"51",
          4427 => x"3f",
          4428 => x"b1",
          4429 => x"3d",
          4430 => x"d6",
          4431 => x"34",
          4432 => x"82",
          4433 => x"a9",
          4434 => x"f6",
          4435 => x"7e",
          4436 => x"72",
          4437 => x"5a",
          4438 => x"2e",
          4439 => x"a2",
          4440 => x"78",
          4441 => x"76",
          4442 => x"81",
          4443 => x"70",
          4444 => x"58",
          4445 => x"2e",
          4446 => x"86",
          4447 => x"26",
          4448 => x"54",
          4449 => x"82",
          4450 => x"70",
          4451 => x"ff",
          4452 => x"82",
          4453 => x"53",
          4454 => x"08",
          4455 => x"f2",
          4456 => x"d8",
          4457 => x"38",
          4458 => x"55",
          4459 => x"88",
          4460 => x"2e",
          4461 => x"39",
          4462 => x"ac",
          4463 => x"5a",
          4464 => x"11",
          4465 => x"51",
          4466 => x"82",
          4467 => x"80",
          4468 => x"ff",
          4469 => x"52",
          4470 => x"b1",
          4471 => x"d8",
          4472 => x"06",
          4473 => x"38",
          4474 => x"39",
          4475 => x"81",
          4476 => x"54",
          4477 => x"ff",
          4478 => x"54",
          4479 => x"d8",
          4480 => x"0d",
          4481 => x"0d",
          4482 => x"b2",
          4483 => x"3d",
          4484 => x"5a",
          4485 => x"3d",
          4486 => x"a4",
          4487 => x"a0",
          4488 => x"73",
          4489 => x"73",
          4490 => x"33",
          4491 => x"83",
          4492 => x"76",
          4493 => x"bc",
          4494 => x"76",
          4495 => x"73",
          4496 => x"ad",
          4497 => x"99",
          4498 => x"d6",
          4499 => x"d5",
          4500 => x"d6",
          4501 => x"2e",
          4502 => x"93",
          4503 => x"82",
          4504 => x"51",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"38",
          4508 => x"51",
          4509 => x"3f",
          4510 => x"82",
          4511 => x"5b",
          4512 => x"08",
          4513 => x"52",
          4514 => x"52",
          4515 => x"a2",
          4516 => x"d8",
          4517 => x"d6",
          4518 => x"2e",
          4519 => x"80",
          4520 => x"d6",
          4521 => x"ff",
          4522 => x"82",
          4523 => x"55",
          4524 => x"d6",
          4525 => x"a9",
          4526 => x"d8",
          4527 => x"70",
          4528 => x"80",
          4529 => x"53",
          4530 => x"06",
          4531 => x"f8",
          4532 => x"1b",
          4533 => x"06",
          4534 => x"7b",
          4535 => x"80",
          4536 => x"2e",
          4537 => x"ff",
          4538 => x"39",
          4539 => x"9c",
          4540 => x"38",
          4541 => x"08",
          4542 => x"38",
          4543 => x"8f",
          4544 => x"c5",
          4545 => x"d8",
          4546 => x"70",
          4547 => x"59",
          4548 => x"ee",
          4549 => x"ff",
          4550 => x"94",
          4551 => x"2b",
          4552 => x"82",
          4553 => x"70",
          4554 => x"97",
          4555 => x"2c",
          4556 => x"29",
          4557 => x"05",
          4558 => x"70",
          4559 => x"51",
          4560 => x"51",
          4561 => x"81",
          4562 => x"2e",
          4563 => x"77",
          4564 => x"38",
          4565 => x"0a",
          4566 => x"0a",
          4567 => x"2c",
          4568 => x"75",
          4569 => x"38",
          4570 => x"52",
          4571 => x"85",
          4572 => x"d8",
          4573 => x"06",
          4574 => x"2e",
          4575 => x"82",
          4576 => x"81",
          4577 => x"74",
          4578 => x"29",
          4579 => x"05",
          4580 => x"70",
          4581 => x"56",
          4582 => x"95",
          4583 => x"76",
          4584 => x"77",
          4585 => x"3f",
          4586 => x"08",
          4587 => x"54",
          4588 => x"d3",
          4589 => x"75",
          4590 => x"ca",
          4591 => x"55",
          4592 => x"94",
          4593 => x"2b",
          4594 => x"82",
          4595 => x"70",
          4596 => x"98",
          4597 => x"11",
          4598 => x"82",
          4599 => x"33",
          4600 => x"51",
          4601 => x"55",
          4602 => x"09",
          4603 => x"92",
          4604 => x"9c",
          4605 => x"0c",
          4606 => x"ee",
          4607 => x"0b",
          4608 => x"34",
          4609 => x"82",
          4610 => x"75",
          4611 => x"34",
          4612 => x"34",
          4613 => x"7e",
          4614 => x"26",
          4615 => x"73",
          4616 => x"ad",
          4617 => x"73",
          4618 => x"ee",
          4619 => x"73",
          4620 => x"cb",
          4621 => x"98",
          4622 => x"75",
          4623 => x"74",
          4624 => x"98",
          4625 => x"73",
          4626 => x"38",
          4627 => x"73",
          4628 => x"34",
          4629 => x"0a",
          4630 => x"0a",
          4631 => x"2c",
          4632 => x"33",
          4633 => x"df",
          4634 => x"9c",
          4635 => x"56",
          4636 => x"ee",
          4637 => x"1a",
          4638 => x"33",
          4639 => x"ee",
          4640 => x"73",
          4641 => x"38",
          4642 => x"73",
          4643 => x"34",
          4644 => x"33",
          4645 => x"0a",
          4646 => x"0a",
          4647 => x"2c",
          4648 => x"33",
          4649 => x"56",
          4650 => x"a8",
          4651 => x"bc",
          4652 => x"1a",
          4653 => x"54",
          4654 => x"3f",
          4655 => x"0a",
          4656 => x"0a",
          4657 => x"2c",
          4658 => x"33",
          4659 => x"73",
          4660 => x"38",
          4661 => x"33",
          4662 => x"70",
          4663 => x"ee",
          4664 => x"51",
          4665 => x"77",
          4666 => x"38",
          4667 => x"08",
          4668 => x"ff",
          4669 => x"74",
          4670 => x"29",
          4671 => x"05",
          4672 => x"82",
          4673 => x"56",
          4674 => x"75",
          4675 => x"fb",
          4676 => x"7a",
          4677 => x"81",
          4678 => x"ee",
          4679 => x"52",
          4680 => x"51",
          4681 => x"81",
          4682 => x"ee",
          4683 => x"81",
          4684 => x"55",
          4685 => x"fb",
          4686 => x"ee",
          4687 => x"05",
          4688 => x"ee",
          4689 => x"15",
          4690 => x"ee",
          4691 => x"f2",
          4692 => x"88",
          4693 => x"da",
          4694 => x"9c",
          4695 => x"2b",
          4696 => x"82",
          4697 => x"57",
          4698 => x"74",
          4699 => x"38",
          4700 => x"81",
          4701 => x"34",
          4702 => x"08",
          4703 => x"51",
          4704 => x"3f",
          4705 => x"0a",
          4706 => x"0a",
          4707 => x"2c",
          4708 => x"33",
          4709 => x"75",
          4710 => x"38",
          4711 => x"08",
          4712 => x"ff",
          4713 => x"82",
          4714 => x"70",
          4715 => x"98",
          4716 => x"98",
          4717 => x"56",
          4718 => x"24",
          4719 => x"82",
          4720 => x"52",
          4721 => x"9f",
          4722 => x"81",
          4723 => x"81",
          4724 => x"70",
          4725 => x"ee",
          4726 => x"51",
          4727 => x"25",
          4728 => x"9b",
          4729 => x"98",
          4730 => x"54",
          4731 => x"82",
          4732 => x"52",
          4733 => x"9f",
          4734 => x"ee",
          4735 => x"51",
          4736 => x"82",
          4737 => x"81",
          4738 => x"73",
          4739 => x"ee",
          4740 => x"73",
          4741 => x"38",
          4742 => x"52",
          4743 => x"f3",
          4744 => x"80",
          4745 => x"0b",
          4746 => x"34",
          4747 => x"ee",
          4748 => x"82",
          4749 => x"af",
          4750 => x"82",
          4751 => x"54",
          4752 => x"f9",
          4753 => x"f2",
          4754 => x"88",
          4755 => x"e2",
          4756 => x"9c",
          4757 => x"54",
          4758 => x"9c",
          4759 => x"ff",
          4760 => x"39",
          4761 => x"33",
          4762 => x"33",
          4763 => x"75",
          4764 => x"38",
          4765 => x"73",
          4766 => x"34",
          4767 => x"70",
          4768 => x"81",
          4769 => x"51",
          4770 => x"25",
          4771 => x"1a",
          4772 => x"33",
          4773 => x"f2",
          4774 => x"73",
          4775 => x"9e",
          4776 => x"81",
          4777 => x"81",
          4778 => x"70",
          4779 => x"ee",
          4780 => x"51",
          4781 => x"24",
          4782 => x"f2",
          4783 => x"a0",
          4784 => x"ee",
          4785 => x"9c",
          4786 => x"2b",
          4787 => x"82",
          4788 => x"57",
          4789 => x"74",
          4790 => x"a3",
          4791 => x"bc",
          4792 => x"51",
          4793 => x"3f",
          4794 => x"0a",
          4795 => x"0a",
          4796 => x"2c",
          4797 => x"33",
          4798 => x"75",
          4799 => x"38",
          4800 => x"82",
          4801 => x"70",
          4802 => x"82",
          4803 => x"59",
          4804 => x"77",
          4805 => x"38",
          4806 => x"08",
          4807 => x"54",
          4808 => x"9c",
          4809 => x"70",
          4810 => x"ff",
          4811 => x"82",
          4812 => x"70",
          4813 => x"82",
          4814 => x"58",
          4815 => x"75",
          4816 => x"f7",
          4817 => x"ee",
          4818 => x"52",
          4819 => x"51",
          4820 => x"80",
          4821 => x"9c",
          4822 => x"82",
          4823 => x"f7",
          4824 => x"b0",
          4825 => x"98",
          4826 => x"80",
          4827 => x"74",
          4828 => x"91",
          4829 => x"d8",
          4830 => x"98",
          4831 => x"d8",
          4832 => x"06",
          4833 => x"74",
          4834 => x"ff",
          4835 => x"93",
          4836 => x"39",
          4837 => x"82",
          4838 => x"fc",
          4839 => x"54",
          4840 => x"a7",
          4841 => x"ff",
          4842 => x"82",
          4843 => x"82",
          4844 => x"82",
          4845 => x"81",
          4846 => x"05",
          4847 => x"79",
          4848 => x"a1",
          4849 => x"54",
          4850 => x"73",
          4851 => x"80",
          4852 => x"38",
          4853 => x"a4",
          4854 => x"39",
          4855 => x"09",
          4856 => x"38",
          4857 => x"08",
          4858 => x"2e",
          4859 => x"51",
          4860 => x"3f",
          4861 => x"08",
          4862 => x"34",
          4863 => x"08",
          4864 => x"81",
          4865 => x"52",
          4866 => x"a5",
          4867 => x"c3",
          4868 => x"29",
          4869 => x"05",
          4870 => x"54",
          4871 => x"ab",
          4872 => x"ff",
          4873 => x"82",
          4874 => x"82",
          4875 => x"82",
          4876 => x"81",
          4877 => x"05",
          4878 => x"79",
          4879 => x"a5",
          4880 => x"54",
          4881 => x"06",
          4882 => x"74",
          4883 => x"34",
          4884 => x"82",
          4885 => x"82",
          4886 => x"52",
          4887 => x"e2",
          4888 => x"39",
          4889 => x"33",
          4890 => x"06",
          4891 => x"33",
          4892 => x"74",
          4893 => x"87",
          4894 => x"bc",
          4895 => x"14",
          4896 => x"ee",
          4897 => x"1a",
          4898 => x"54",
          4899 => x"3f",
          4900 => x"82",
          4901 => x"54",
          4902 => x"f4",
          4903 => x"f2",
          4904 => x"88",
          4905 => x"8a",
          4906 => x"9c",
          4907 => x"54",
          4908 => x"9c",
          4909 => x"39",
          4910 => x"02",
          4911 => x"52",
          4912 => x"09",
          4913 => x"38",
          4914 => x"08",
          4915 => x"d6",
          4916 => x"0b",
          4917 => x"08",
          4918 => x"98",
          4919 => x"c4",
          4920 => x"82",
          4921 => x"82",
          4922 => x"84",
          4923 => x"c4",
          4924 => x"88",
          4925 => x"c8",
          4926 => x"a0",
          4927 => x"70",
          4928 => x"0c",
          4929 => x"82",
          4930 => x"33",
          4931 => x"d6",
          4932 => x"05",
          4933 => x"0c",
          4934 => x"d6",
          4935 => x"a0",
          4936 => x"c4",
          4937 => x"82",
          4938 => x"98",
          4939 => x"c4",
          4940 => x"38",
          4941 => x"d6",
          4942 => x"0b",
          4943 => x"0c",
          4944 => x"d6",
          4945 => x"3d",
          4946 => x"0b",
          4947 => x"0c",
          4948 => x"0d",
          4949 => x"0b",
          4950 => x"0c",
          4951 => x"82",
          4952 => x"a0",
          4953 => x"52",
          4954 => x"51",
          4955 => x"3f",
          4956 => x"08",
          4957 => x"77",
          4958 => x"57",
          4959 => x"34",
          4960 => x"08",
          4961 => x"15",
          4962 => x"15",
          4963 => x"d0",
          4964 => x"86",
          4965 => x"87",
          4966 => x"d6",
          4967 => x"d6",
          4968 => x"05",
          4969 => x"07",
          4970 => x"ff",
          4971 => x"2a",
          4972 => x"56",
          4973 => x"34",
          4974 => x"34",
          4975 => x"22",
          4976 => x"82",
          4977 => x"05",
          4978 => x"55",
          4979 => x"15",
          4980 => x"15",
          4981 => x"0d",
          4982 => x"0d",
          4983 => x"51",
          4984 => x"8f",
          4985 => x"83",
          4986 => x"70",
          4987 => x"06",
          4988 => x"70",
          4989 => x"0c",
          4990 => x"04",
          4991 => x"02",
          4992 => x"02",
          4993 => x"05",
          4994 => x"82",
          4995 => x"71",
          4996 => x"11",
          4997 => x"73",
          4998 => x"81",
          4999 => x"88",
          5000 => x"a4",
          5001 => x"22",
          5002 => x"ff",
          5003 => x"88",
          5004 => x"52",
          5005 => x"5b",
          5006 => x"55",
          5007 => x"70",
          5008 => x"82",
          5009 => x"14",
          5010 => x"52",
          5011 => x"15",
          5012 => x"15",
          5013 => x"d0",
          5014 => x"70",
          5015 => x"33",
          5016 => x"07",
          5017 => x"8f",
          5018 => x"51",
          5019 => x"71",
          5020 => x"ff",
          5021 => x"88",
          5022 => x"51",
          5023 => x"34",
          5024 => x"06",
          5025 => x"12",
          5026 => x"d0",
          5027 => x"71",
          5028 => x"81",
          5029 => x"3d",
          5030 => x"3d",
          5031 => x"d0",
          5032 => x"05",
          5033 => x"70",
          5034 => x"11",
          5035 => x"87",
          5036 => x"8b",
          5037 => x"2b",
          5038 => x"59",
          5039 => x"72",
          5040 => x"33",
          5041 => x"71",
          5042 => x"70",
          5043 => x"56",
          5044 => x"84",
          5045 => x"85",
          5046 => x"d6",
          5047 => x"14",
          5048 => x"85",
          5049 => x"8b",
          5050 => x"2b",
          5051 => x"57",
          5052 => x"86",
          5053 => x"13",
          5054 => x"2b",
          5055 => x"2a",
          5056 => x"52",
          5057 => x"34",
          5058 => x"34",
          5059 => x"08",
          5060 => x"81",
          5061 => x"88",
          5062 => x"81",
          5063 => x"70",
          5064 => x"51",
          5065 => x"71",
          5066 => x"81",
          5067 => x"3d",
          5068 => x"3d",
          5069 => x"05",
          5070 => x"d0",
          5071 => x"2b",
          5072 => x"33",
          5073 => x"71",
          5074 => x"70",
          5075 => x"70",
          5076 => x"33",
          5077 => x"71",
          5078 => x"53",
          5079 => x"52",
          5080 => x"53",
          5081 => x"25",
          5082 => x"72",
          5083 => x"3f",
          5084 => x"08",
          5085 => x"33",
          5086 => x"71",
          5087 => x"83",
          5088 => x"11",
          5089 => x"12",
          5090 => x"2b",
          5091 => x"2b",
          5092 => x"06",
          5093 => x"51",
          5094 => x"53",
          5095 => x"88",
          5096 => x"72",
          5097 => x"73",
          5098 => x"82",
          5099 => x"70",
          5100 => x"81",
          5101 => x"8b",
          5102 => x"2b",
          5103 => x"57",
          5104 => x"70",
          5105 => x"33",
          5106 => x"07",
          5107 => x"ff",
          5108 => x"2a",
          5109 => x"58",
          5110 => x"34",
          5111 => x"34",
          5112 => x"04",
          5113 => x"82",
          5114 => x"02",
          5115 => x"05",
          5116 => x"2b",
          5117 => x"11",
          5118 => x"33",
          5119 => x"71",
          5120 => x"59",
          5121 => x"56",
          5122 => x"71",
          5123 => x"33",
          5124 => x"07",
          5125 => x"a2",
          5126 => x"07",
          5127 => x"53",
          5128 => x"53",
          5129 => x"70",
          5130 => x"82",
          5131 => x"70",
          5132 => x"81",
          5133 => x"8b",
          5134 => x"2b",
          5135 => x"57",
          5136 => x"82",
          5137 => x"13",
          5138 => x"2b",
          5139 => x"2a",
          5140 => x"52",
          5141 => x"34",
          5142 => x"34",
          5143 => x"08",
          5144 => x"33",
          5145 => x"71",
          5146 => x"82",
          5147 => x"52",
          5148 => x"0d",
          5149 => x"0d",
          5150 => x"d0",
          5151 => x"2a",
          5152 => x"ff",
          5153 => x"57",
          5154 => x"3f",
          5155 => x"08",
          5156 => x"71",
          5157 => x"33",
          5158 => x"71",
          5159 => x"83",
          5160 => x"11",
          5161 => x"12",
          5162 => x"2b",
          5163 => x"07",
          5164 => x"51",
          5165 => x"55",
          5166 => x"80",
          5167 => x"82",
          5168 => x"75",
          5169 => x"3f",
          5170 => x"84",
          5171 => x"15",
          5172 => x"2b",
          5173 => x"07",
          5174 => x"88",
          5175 => x"55",
          5176 => x"86",
          5177 => x"81",
          5178 => x"75",
          5179 => x"82",
          5180 => x"70",
          5181 => x"33",
          5182 => x"71",
          5183 => x"70",
          5184 => x"57",
          5185 => x"72",
          5186 => x"73",
          5187 => x"82",
          5188 => x"18",
          5189 => x"86",
          5190 => x"0b",
          5191 => x"82",
          5192 => x"53",
          5193 => x"34",
          5194 => x"34",
          5195 => x"08",
          5196 => x"81",
          5197 => x"88",
          5198 => x"82",
          5199 => x"70",
          5200 => x"51",
          5201 => x"74",
          5202 => x"81",
          5203 => x"3d",
          5204 => x"3d",
          5205 => x"82",
          5206 => x"84",
          5207 => x"3f",
          5208 => x"86",
          5209 => x"fe",
          5210 => x"3d",
          5211 => x"3d",
          5212 => x"52",
          5213 => x"3f",
          5214 => x"08",
          5215 => x"06",
          5216 => x"08",
          5217 => x"85",
          5218 => x"88",
          5219 => x"5f",
          5220 => x"5a",
          5221 => x"59",
          5222 => x"80",
          5223 => x"88",
          5224 => x"33",
          5225 => x"71",
          5226 => x"70",
          5227 => x"06",
          5228 => x"83",
          5229 => x"70",
          5230 => x"53",
          5231 => x"55",
          5232 => x"8a",
          5233 => x"2e",
          5234 => x"78",
          5235 => x"15",
          5236 => x"33",
          5237 => x"07",
          5238 => x"c2",
          5239 => x"ff",
          5240 => x"38",
          5241 => x"56",
          5242 => x"2b",
          5243 => x"08",
          5244 => x"81",
          5245 => x"88",
          5246 => x"81",
          5247 => x"51",
          5248 => x"5c",
          5249 => x"2e",
          5250 => x"55",
          5251 => x"78",
          5252 => x"38",
          5253 => x"80",
          5254 => x"38",
          5255 => x"09",
          5256 => x"38",
          5257 => x"f2",
          5258 => x"39",
          5259 => x"53",
          5260 => x"51",
          5261 => x"82",
          5262 => x"70",
          5263 => x"33",
          5264 => x"71",
          5265 => x"83",
          5266 => x"5a",
          5267 => x"05",
          5268 => x"83",
          5269 => x"70",
          5270 => x"59",
          5271 => x"84",
          5272 => x"81",
          5273 => x"76",
          5274 => x"82",
          5275 => x"75",
          5276 => x"11",
          5277 => x"11",
          5278 => x"33",
          5279 => x"07",
          5280 => x"53",
          5281 => x"5a",
          5282 => x"86",
          5283 => x"87",
          5284 => x"d6",
          5285 => x"1c",
          5286 => x"85",
          5287 => x"8b",
          5288 => x"2b",
          5289 => x"5a",
          5290 => x"54",
          5291 => x"34",
          5292 => x"34",
          5293 => x"08",
          5294 => x"1d",
          5295 => x"85",
          5296 => x"88",
          5297 => x"88",
          5298 => x"5f",
          5299 => x"73",
          5300 => x"75",
          5301 => x"82",
          5302 => x"1b",
          5303 => x"73",
          5304 => x"0c",
          5305 => x"04",
          5306 => x"74",
          5307 => x"d0",
          5308 => x"f4",
          5309 => x"53",
          5310 => x"8b",
          5311 => x"fc",
          5312 => x"d6",
          5313 => x"72",
          5314 => x"0c",
          5315 => x"04",
          5316 => x"64",
          5317 => x"80",
          5318 => x"82",
          5319 => x"60",
          5320 => x"06",
          5321 => x"a9",
          5322 => x"38",
          5323 => x"b8",
          5324 => x"d8",
          5325 => x"c7",
          5326 => x"38",
          5327 => x"92",
          5328 => x"83",
          5329 => x"51",
          5330 => x"82",
          5331 => x"83",
          5332 => x"82",
          5333 => x"7d",
          5334 => x"2a",
          5335 => x"ff",
          5336 => x"2b",
          5337 => x"33",
          5338 => x"71",
          5339 => x"70",
          5340 => x"83",
          5341 => x"70",
          5342 => x"05",
          5343 => x"1a",
          5344 => x"12",
          5345 => x"2b",
          5346 => x"2b",
          5347 => x"53",
          5348 => x"5c",
          5349 => x"5c",
          5350 => x"73",
          5351 => x"38",
          5352 => x"ff",
          5353 => x"70",
          5354 => x"06",
          5355 => x"16",
          5356 => x"33",
          5357 => x"07",
          5358 => x"1c",
          5359 => x"12",
          5360 => x"2b",
          5361 => x"07",
          5362 => x"52",
          5363 => x"80",
          5364 => x"78",
          5365 => x"83",
          5366 => x"41",
          5367 => x"27",
          5368 => x"60",
          5369 => x"7b",
          5370 => x"06",
          5371 => x"51",
          5372 => x"7a",
          5373 => x"06",
          5374 => x"39",
          5375 => x"7a",
          5376 => x"38",
          5377 => x"aa",
          5378 => x"39",
          5379 => x"7a",
          5380 => x"c8",
          5381 => x"82",
          5382 => x"12",
          5383 => x"2b",
          5384 => x"54",
          5385 => x"80",
          5386 => x"f7",
          5387 => x"d6",
          5388 => x"ff",
          5389 => x"54",
          5390 => x"83",
          5391 => x"d0",
          5392 => x"05",
          5393 => x"ff",
          5394 => x"82",
          5395 => x"14",
          5396 => x"83",
          5397 => x"59",
          5398 => x"39",
          5399 => x"7a",
          5400 => x"d4",
          5401 => x"f5",
          5402 => x"d6",
          5403 => x"82",
          5404 => x"12",
          5405 => x"2b",
          5406 => x"54",
          5407 => x"80",
          5408 => x"f6",
          5409 => x"d6",
          5410 => x"ff",
          5411 => x"54",
          5412 => x"83",
          5413 => x"d0",
          5414 => x"05",
          5415 => x"ff",
          5416 => x"82",
          5417 => x"14",
          5418 => x"62",
          5419 => x"5c",
          5420 => x"ff",
          5421 => x"39",
          5422 => x"54",
          5423 => x"82",
          5424 => x"5c",
          5425 => x"08",
          5426 => x"38",
          5427 => x"52",
          5428 => x"08",
          5429 => x"8d",
          5430 => x"f7",
          5431 => x"58",
          5432 => x"99",
          5433 => x"7a",
          5434 => x"f2",
          5435 => x"19",
          5436 => x"d6",
          5437 => x"84",
          5438 => x"f9",
          5439 => x"73",
          5440 => x"0c",
          5441 => x"04",
          5442 => x"77",
          5443 => x"52",
          5444 => x"3f",
          5445 => x"08",
          5446 => x"d8",
          5447 => x"8e",
          5448 => x"80",
          5449 => x"d8",
          5450 => x"99",
          5451 => x"82",
          5452 => x"86",
          5453 => x"ff",
          5454 => x"8f",
          5455 => x"81",
          5456 => x"26",
          5457 => x"d6",
          5458 => x"52",
          5459 => x"d8",
          5460 => x"0d",
          5461 => x"0d",
          5462 => x"33",
          5463 => x"9f",
          5464 => x"53",
          5465 => x"81",
          5466 => x"38",
          5467 => x"87",
          5468 => x"11",
          5469 => x"54",
          5470 => x"84",
          5471 => x"54",
          5472 => x"87",
          5473 => x"11",
          5474 => x"0c",
          5475 => x"c0",
          5476 => x"70",
          5477 => x"70",
          5478 => x"51",
          5479 => x"8a",
          5480 => x"98",
          5481 => x"70",
          5482 => x"08",
          5483 => x"06",
          5484 => x"38",
          5485 => x"8c",
          5486 => x"80",
          5487 => x"71",
          5488 => x"14",
          5489 => x"d4",
          5490 => x"70",
          5491 => x"0c",
          5492 => x"04",
          5493 => x"60",
          5494 => x"8c",
          5495 => x"33",
          5496 => x"5b",
          5497 => x"5a",
          5498 => x"82",
          5499 => x"81",
          5500 => x"52",
          5501 => x"38",
          5502 => x"84",
          5503 => x"92",
          5504 => x"c0",
          5505 => x"87",
          5506 => x"13",
          5507 => x"57",
          5508 => x"0b",
          5509 => x"8c",
          5510 => x"0c",
          5511 => x"75",
          5512 => x"2a",
          5513 => x"51",
          5514 => x"80",
          5515 => x"7b",
          5516 => x"7b",
          5517 => x"5d",
          5518 => x"59",
          5519 => x"06",
          5520 => x"73",
          5521 => x"81",
          5522 => x"ff",
          5523 => x"72",
          5524 => x"38",
          5525 => x"8c",
          5526 => x"c3",
          5527 => x"98",
          5528 => x"71",
          5529 => x"38",
          5530 => x"2e",
          5531 => x"76",
          5532 => x"92",
          5533 => x"72",
          5534 => x"06",
          5535 => x"f7",
          5536 => x"5a",
          5537 => x"80",
          5538 => x"70",
          5539 => x"5a",
          5540 => x"80",
          5541 => x"73",
          5542 => x"06",
          5543 => x"38",
          5544 => x"fe",
          5545 => x"fc",
          5546 => x"52",
          5547 => x"83",
          5548 => x"71",
          5549 => x"d6",
          5550 => x"3d",
          5551 => x"3d",
          5552 => x"64",
          5553 => x"bf",
          5554 => x"40",
          5555 => x"59",
          5556 => x"58",
          5557 => x"82",
          5558 => x"81",
          5559 => x"52",
          5560 => x"09",
          5561 => x"b1",
          5562 => x"84",
          5563 => x"92",
          5564 => x"c0",
          5565 => x"87",
          5566 => x"13",
          5567 => x"56",
          5568 => x"87",
          5569 => x"0c",
          5570 => x"82",
          5571 => x"58",
          5572 => x"84",
          5573 => x"06",
          5574 => x"71",
          5575 => x"38",
          5576 => x"05",
          5577 => x"0c",
          5578 => x"73",
          5579 => x"81",
          5580 => x"71",
          5581 => x"38",
          5582 => x"8c",
          5583 => x"d0",
          5584 => x"98",
          5585 => x"71",
          5586 => x"38",
          5587 => x"2e",
          5588 => x"76",
          5589 => x"92",
          5590 => x"72",
          5591 => x"06",
          5592 => x"f7",
          5593 => x"59",
          5594 => x"1a",
          5595 => x"06",
          5596 => x"59",
          5597 => x"80",
          5598 => x"73",
          5599 => x"06",
          5600 => x"38",
          5601 => x"fe",
          5602 => x"fc",
          5603 => x"52",
          5604 => x"83",
          5605 => x"71",
          5606 => x"d6",
          5607 => x"3d",
          5608 => x"3d",
          5609 => x"84",
          5610 => x"33",
          5611 => x"a7",
          5612 => x"54",
          5613 => x"fa",
          5614 => x"d6",
          5615 => x"06",
          5616 => x"72",
          5617 => x"85",
          5618 => x"98",
          5619 => x"56",
          5620 => x"80",
          5621 => x"76",
          5622 => x"74",
          5623 => x"c0",
          5624 => x"54",
          5625 => x"2e",
          5626 => x"d4",
          5627 => x"2e",
          5628 => x"80",
          5629 => x"08",
          5630 => x"70",
          5631 => x"51",
          5632 => x"2e",
          5633 => x"c0",
          5634 => x"52",
          5635 => x"87",
          5636 => x"08",
          5637 => x"38",
          5638 => x"87",
          5639 => x"14",
          5640 => x"70",
          5641 => x"52",
          5642 => x"96",
          5643 => x"92",
          5644 => x"0a",
          5645 => x"39",
          5646 => x"0c",
          5647 => x"39",
          5648 => x"54",
          5649 => x"d8",
          5650 => x"0d",
          5651 => x"0d",
          5652 => x"33",
          5653 => x"88",
          5654 => x"d6",
          5655 => x"51",
          5656 => x"04",
          5657 => x"75",
          5658 => x"82",
          5659 => x"90",
          5660 => x"2b",
          5661 => x"33",
          5662 => x"88",
          5663 => x"71",
          5664 => x"d8",
          5665 => x"54",
          5666 => x"85",
          5667 => x"ff",
          5668 => x"02",
          5669 => x"05",
          5670 => x"70",
          5671 => x"05",
          5672 => x"88",
          5673 => x"72",
          5674 => x"0d",
          5675 => x"0d",
          5676 => x"52",
          5677 => x"81",
          5678 => x"70",
          5679 => x"70",
          5680 => x"05",
          5681 => x"88",
          5682 => x"72",
          5683 => x"54",
          5684 => x"2a",
          5685 => x"34",
          5686 => x"04",
          5687 => x"76",
          5688 => x"54",
          5689 => x"2e",
          5690 => x"70",
          5691 => x"33",
          5692 => x"05",
          5693 => x"11",
          5694 => x"84",
          5695 => x"fe",
          5696 => x"77",
          5697 => x"53",
          5698 => x"81",
          5699 => x"ff",
          5700 => x"f4",
          5701 => x"0d",
          5702 => x"0d",
          5703 => x"56",
          5704 => x"70",
          5705 => x"33",
          5706 => x"05",
          5707 => x"71",
          5708 => x"56",
          5709 => x"72",
          5710 => x"38",
          5711 => x"e2",
          5712 => x"d6",
          5713 => x"3d",
          5714 => x"3d",
          5715 => x"54",
          5716 => x"71",
          5717 => x"38",
          5718 => x"70",
          5719 => x"f3",
          5720 => x"82",
          5721 => x"84",
          5722 => x"80",
          5723 => x"d8",
          5724 => x"3d",
          5725 => x"08",
          5726 => x"05",
          5727 => x"54",
          5728 => x"e7",
          5729 => x"82",
          5730 => x"a2",
          5731 => x"2e",
          5732 => x"b5",
          5733 => x"80",
          5734 => x"82",
          5735 => x"83",
          5736 => x"53",
          5737 => x"86",
          5738 => x"0c",
          5739 => x"82",
          5740 => x"87",
          5741 => x"f7",
          5742 => x"56",
          5743 => x"17",
          5744 => x"74",
          5745 => x"d6",
          5746 => x"b4",
          5747 => x"b8",
          5748 => x"81",
          5749 => x"59",
          5750 => x"82",
          5751 => x"7a",
          5752 => x"06",
          5753 => x"d6",
          5754 => x"17",
          5755 => x"08",
          5756 => x"08",
          5757 => x"08",
          5758 => x"74",
          5759 => x"38",
          5760 => x"55",
          5761 => x"09",
          5762 => x"38",
          5763 => x"18",
          5764 => x"81",
          5765 => x"f9",
          5766 => x"39",
          5767 => x"82",
          5768 => x"8b",
          5769 => x"fa",
          5770 => x"7a",
          5771 => x"57",
          5772 => x"08",
          5773 => x"75",
          5774 => x"3f",
          5775 => x"08",
          5776 => x"d8",
          5777 => x"81",
          5778 => x"b8",
          5779 => x"16",
          5780 => x"80",
          5781 => x"d8",
          5782 => x"85",
          5783 => x"81",
          5784 => x"17",
          5785 => x"d6",
          5786 => x"3d",
          5787 => x"3d",
          5788 => x"52",
          5789 => x"3f",
          5790 => x"08",
          5791 => x"d8",
          5792 => x"38",
          5793 => x"74",
          5794 => x"81",
          5795 => x"38",
          5796 => x"59",
          5797 => x"09",
          5798 => x"e3",
          5799 => x"53",
          5800 => x"08",
          5801 => x"70",
          5802 => x"d3",
          5803 => x"d5",
          5804 => x"17",
          5805 => x"3f",
          5806 => x"a4",
          5807 => x"51",
          5808 => x"86",
          5809 => x"f2",
          5810 => x"17",
          5811 => x"3f",
          5812 => x"52",
          5813 => x"51",
          5814 => x"90",
          5815 => x"84",
          5816 => x"fb",
          5817 => x"17",
          5818 => x"70",
          5819 => x"79",
          5820 => x"52",
          5821 => x"51",
          5822 => x"77",
          5823 => x"80",
          5824 => x"81",
          5825 => x"f9",
          5826 => x"d6",
          5827 => x"2e",
          5828 => x"58",
          5829 => x"d8",
          5830 => x"0d",
          5831 => x"0d",
          5832 => x"9c",
          5833 => x"05",
          5834 => x"80",
          5835 => x"27",
          5836 => x"14",
          5837 => x"29",
          5838 => x"05",
          5839 => x"82",
          5840 => x"87",
          5841 => x"f9",
          5842 => x"7a",
          5843 => x"54",
          5844 => x"27",
          5845 => x"76",
          5846 => x"27",
          5847 => x"ff",
          5848 => x"58",
          5849 => x"80",
          5850 => x"82",
          5851 => x"72",
          5852 => x"38",
          5853 => x"72",
          5854 => x"8e",
          5855 => x"39",
          5856 => x"17",
          5857 => x"a8",
          5858 => x"53",
          5859 => x"fd",
          5860 => x"d6",
          5861 => x"9f",
          5862 => x"ff",
          5863 => x"11",
          5864 => x"70",
          5865 => x"18",
          5866 => x"76",
          5867 => x"53",
          5868 => x"82",
          5869 => x"80",
          5870 => x"83",
          5871 => x"b8",
          5872 => x"88",
          5873 => x"79",
          5874 => x"84",
          5875 => x"58",
          5876 => x"80",
          5877 => x"9f",
          5878 => x"80",
          5879 => x"88",
          5880 => x"08",
          5881 => x"51",
          5882 => x"82",
          5883 => x"80",
          5884 => x"10",
          5885 => x"74",
          5886 => x"51",
          5887 => x"82",
          5888 => x"83",
          5889 => x"58",
          5890 => x"87",
          5891 => x"08",
          5892 => x"51",
          5893 => x"82",
          5894 => x"9b",
          5895 => x"2b",
          5896 => x"74",
          5897 => x"51",
          5898 => x"82",
          5899 => x"f0",
          5900 => x"83",
          5901 => x"77",
          5902 => x"0c",
          5903 => x"04",
          5904 => x"7a",
          5905 => x"58",
          5906 => x"81",
          5907 => x"9e",
          5908 => x"17",
          5909 => x"96",
          5910 => x"53",
          5911 => x"81",
          5912 => x"79",
          5913 => x"72",
          5914 => x"38",
          5915 => x"72",
          5916 => x"b8",
          5917 => x"39",
          5918 => x"17",
          5919 => x"a8",
          5920 => x"53",
          5921 => x"fb",
          5922 => x"d6",
          5923 => x"82",
          5924 => x"81",
          5925 => x"83",
          5926 => x"b8",
          5927 => x"78",
          5928 => x"56",
          5929 => x"76",
          5930 => x"38",
          5931 => x"9f",
          5932 => x"33",
          5933 => x"07",
          5934 => x"74",
          5935 => x"83",
          5936 => x"89",
          5937 => x"08",
          5938 => x"51",
          5939 => x"82",
          5940 => x"59",
          5941 => x"08",
          5942 => x"74",
          5943 => x"16",
          5944 => x"84",
          5945 => x"76",
          5946 => x"88",
          5947 => x"81",
          5948 => x"8f",
          5949 => x"53",
          5950 => x"80",
          5951 => x"88",
          5952 => x"08",
          5953 => x"51",
          5954 => x"82",
          5955 => x"59",
          5956 => x"08",
          5957 => x"77",
          5958 => x"06",
          5959 => x"83",
          5960 => x"05",
          5961 => x"f6",
          5962 => x"39",
          5963 => x"a8",
          5964 => x"52",
          5965 => x"ef",
          5966 => x"d8",
          5967 => x"d6",
          5968 => x"38",
          5969 => x"06",
          5970 => x"83",
          5971 => x"18",
          5972 => x"54",
          5973 => x"f6",
          5974 => x"d6",
          5975 => x"0a",
          5976 => x"52",
          5977 => x"c5",
          5978 => x"83",
          5979 => x"82",
          5980 => x"8a",
          5981 => x"f8",
          5982 => x"7c",
          5983 => x"59",
          5984 => x"81",
          5985 => x"38",
          5986 => x"08",
          5987 => x"73",
          5988 => x"38",
          5989 => x"52",
          5990 => x"a4",
          5991 => x"d8",
          5992 => x"d6",
          5993 => x"f2",
          5994 => x"82",
          5995 => x"39",
          5996 => x"e6",
          5997 => x"d8",
          5998 => x"de",
          5999 => x"78",
          6000 => x"3f",
          6001 => x"08",
          6002 => x"d8",
          6003 => x"80",
          6004 => x"d6",
          6005 => x"2e",
          6006 => x"d6",
          6007 => x"2e",
          6008 => x"53",
          6009 => x"51",
          6010 => x"82",
          6011 => x"c5",
          6012 => x"08",
          6013 => x"18",
          6014 => x"57",
          6015 => x"90",
          6016 => x"94",
          6017 => x"16",
          6018 => x"54",
          6019 => x"34",
          6020 => x"78",
          6021 => x"38",
          6022 => x"82",
          6023 => x"8a",
          6024 => x"f6",
          6025 => x"7e",
          6026 => x"5b",
          6027 => x"38",
          6028 => x"58",
          6029 => x"88",
          6030 => x"08",
          6031 => x"38",
          6032 => x"39",
          6033 => x"51",
          6034 => x"81",
          6035 => x"d6",
          6036 => x"82",
          6037 => x"d6",
          6038 => x"82",
          6039 => x"ff",
          6040 => x"38",
          6041 => x"82",
          6042 => x"26",
          6043 => x"79",
          6044 => x"08",
          6045 => x"73",
          6046 => x"b9",
          6047 => x"2e",
          6048 => x"80",
          6049 => x"1a",
          6050 => x"08",
          6051 => x"38",
          6052 => x"52",
          6053 => x"af",
          6054 => x"82",
          6055 => x"81",
          6056 => x"06",
          6057 => x"d6",
          6058 => x"82",
          6059 => x"09",
          6060 => x"72",
          6061 => x"70",
          6062 => x"d6",
          6063 => x"51",
          6064 => x"73",
          6065 => x"82",
          6066 => x"80",
          6067 => x"90",
          6068 => x"81",
          6069 => x"38",
          6070 => x"08",
          6071 => x"73",
          6072 => x"75",
          6073 => x"77",
          6074 => x"56",
          6075 => x"76",
          6076 => x"82",
          6077 => x"26",
          6078 => x"75",
          6079 => x"f8",
          6080 => x"d6",
          6081 => x"2e",
          6082 => x"59",
          6083 => x"08",
          6084 => x"81",
          6085 => x"82",
          6086 => x"59",
          6087 => x"08",
          6088 => x"70",
          6089 => x"25",
          6090 => x"51",
          6091 => x"73",
          6092 => x"75",
          6093 => x"81",
          6094 => x"38",
          6095 => x"f5",
          6096 => x"75",
          6097 => x"f9",
          6098 => x"d6",
          6099 => x"d6",
          6100 => x"70",
          6101 => x"08",
          6102 => x"51",
          6103 => x"80",
          6104 => x"73",
          6105 => x"38",
          6106 => x"52",
          6107 => x"d0",
          6108 => x"d8",
          6109 => x"a5",
          6110 => x"18",
          6111 => x"08",
          6112 => x"18",
          6113 => x"74",
          6114 => x"38",
          6115 => x"18",
          6116 => x"33",
          6117 => x"73",
          6118 => x"97",
          6119 => x"74",
          6120 => x"38",
          6121 => x"55",
          6122 => x"d6",
          6123 => x"85",
          6124 => x"75",
          6125 => x"d6",
          6126 => x"3d",
          6127 => x"3d",
          6128 => x"52",
          6129 => x"3f",
          6130 => x"08",
          6131 => x"82",
          6132 => x"80",
          6133 => x"52",
          6134 => x"c1",
          6135 => x"d8",
          6136 => x"d8",
          6137 => x"0c",
          6138 => x"53",
          6139 => x"15",
          6140 => x"f2",
          6141 => x"56",
          6142 => x"16",
          6143 => x"22",
          6144 => x"27",
          6145 => x"54",
          6146 => x"76",
          6147 => x"33",
          6148 => x"3f",
          6149 => x"08",
          6150 => x"38",
          6151 => x"76",
          6152 => x"70",
          6153 => x"9f",
          6154 => x"56",
          6155 => x"d6",
          6156 => x"3d",
          6157 => x"3d",
          6158 => x"71",
          6159 => x"57",
          6160 => x"0a",
          6161 => x"38",
          6162 => x"53",
          6163 => x"38",
          6164 => x"0c",
          6165 => x"54",
          6166 => x"75",
          6167 => x"73",
          6168 => x"ac",
          6169 => x"73",
          6170 => x"85",
          6171 => x"0b",
          6172 => x"5a",
          6173 => x"27",
          6174 => x"ac",
          6175 => x"18",
          6176 => x"39",
          6177 => x"70",
          6178 => x"58",
          6179 => x"b2",
          6180 => x"76",
          6181 => x"3f",
          6182 => x"08",
          6183 => x"d8",
          6184 => x"bd",
          6185 => x"82",
          6186 => x"27",
          6187 => x"16",
          6188 => x"d8",
          6189 => x"38",
          6190 => x"39",
          6191 => x"55",
          6192 => x"52",
          6193 => x"d5",
          6194 => x"d8",
          6195 => x"0c",
          6196 => x"0c",
          6197 => x"53",
          6198 => x"80",
          6199 => x"85",
          6200 => x"94",
          6201 => x"2a",
          6202 => x"0c",
          6203 => x"06",
          6204 => x"9c",
          6205 => x"58",
          6206 => x"d8",
          6207 => x"0d",
          6208 => x"0d",
          6209 => x"90",
          6210 => x"05",
          6211 => x"f0",
          6212 => x"27",
          6213 => x"0b",
          6214 => x"98",
          6215 => x"84",
          6216 => x"2e",
          6217 => x"76",
          6218 => x"58",
          6219 => x"38",
          6220 => x"15",
          6221 => x"08",
          6222 => x"38",
          6223 => x"88",
          6224 => x"53",
          6225 => x"81",
          6226 => x"c0",
          6227 => x"22",
          6228 => x"89",
          6229 => x"72",
          6230 => x"74",
          6231 => x"f3",
          6232 => x"d6",
          6233 => x"82",
          6234 => x"82",
          6235 => x"27",
          6236 => x"81",
          6237 => x"d8",
          6238 => x"80",
          6239 => x"16",
          6240 => x"d8",
          6241 => x"ca",
          6242 => x"38",
          6243 => x"0c",
          6244 => x"dd",
          6245 => x"08",
          6246 => x"f9",
          6247 => x"d6",
          6248 => x"87",
          6249 => x"d8",
          6250 => x"80",
          6251 => x"55",
          6252 => x"08",
          6253 => x"38",
          6254 => x"d6",
          6255 => x"2e",
          6256 => x"d6",
          6257 => x"75",
          6258 => x"3f",
          6259 => x"08",
          6260 => x"94",
          6261 => x"52",
          6262 => x"c1",
          6263 => x"d8",
          6264 => x"0c",
          6265 => x"0c",
          6266 => x"05",
          6267 => x"80",
          6268 => x"d6",
          6269 => x"3d",
          6270 => x"3d",
          6271 => x"71",
          6272 => x"57",
          6273 => x"51",
          6274 => x"82",
          6275 => x"54",
          6276 => x"08",
          6277 => x"82",
          6278 => x"56",
          6279 => x"52",
          6280 => x"83",
          6281 => x"d8",
          6282 => x"d6",
          6283 => x"d2",
          6284 => x"d8",
          6285 => x"08",
          6286 => x"54",
          6287 => x"e5",
          6288 => x"06",
          6289 => x"58",
          6290 => x"08",
          6291 => x"38",
          6292 => x"75",
          6293 => x"80",
          6294 => x"81",
          6295 => x"7a",
          6296 => x"06",
          6297 => x"39",
          6298 => x"08",
          6299 => x"76",
          6300 => x"3f",
          6301 => x"08",
          6302 => x"d8",
          6303 => x"ff",
          6304 => x"84",
          6305 => x"06",
          6306 => x"54",
          6307 => x"d8",
          6308 => x"0d",
          6309 => x"0d",
          6310 => x"52",
          6311 => x"3f",
          6312 => x"08",
          6313 => x"06",
          6314 => x"51",
          6315 => x"83",
          6316 => x"06",
          6317 => x"14",
          6318 => x"3f",
          6319 => x"08",
          6320 => x"07",
          6321 => x"d6",
          6322 => x"3d",
          6323 => x"3d",
          6324 => x"70",
          6325 => x"06",
          6326 => x"53",
          6327 => x"af",
          6328 => x"33",
          6329 => x"83",
          6330 => x"06",
          6331 => x"90",
          6332 => x"15",
          6333 => x"3f",
          6334 => x"04",
          6335 => x"75",
          6336 => x"8b",
          6337 => x"2a",
          6338 => x"29",
          6339 => x"81",
          6340 => x"71",
          6341 => x"ff",
          6342 => x"56",
          6343 => x"72",
          6344 => x"82",
          6345 => x"85",
          6346 => x"f2",
          6347 => x"62",
          6348 => x"79",
          6349 => x"81",
          6350 => x"5d",
          6351 => x"80",
          6352 => x"38",
          6353 => x"52",
          6354 => x"db",
          6355 => x"d8",
          6356 => x"d6",
          6357 => x"eb",
          6358 => x"08",
          6359 => x"55",
          6360 => x"84",
          6361 => x"39",
          6362 => x"bf",
          6363 => x"ff",
          6364 => x"72",
          6365 => x"82",
          6366 => x"56",
          6367 => x"2e",
          6368 => x"83",
          6369 => x"82",
          6370 => x"53",
          6371 => x"09",
          6372 => x"38",
          6373 => x"73",
          6374 => x"99",
          6375 => x"d8",
          6376 => x"06",
          6377 => x"88",
          6378 => x"06",
          6379 => x"56",
          6380 => x"87",
          6381 => x"5c",
          6382 => x"76",
          6383 => x"81",
          6384 => x"38",
          6385 => x"70",
          6386 => x"53",
          6387 => x"92",
          6388 => x"33",
          6389 => x"06",
          6390 => x"08",
          6391 => x"56",
          6392 => x"7c",
          6393 => x"06",
          6394 => x"8d",
          6395 => x"7c",
          6396 => x"81",
          6397 => x"38",
          6398 => x"9a",
          6399 => x"e8",
          6400 => x"d6",
          6401 => x"ff",
          6402 => x"72",
          6403 => x"74",
          6404 => x"bf",
          6405 => x"f3",
          6406 => x"81",
          6407 => x"82",
          6408 => x"33",
          6409 => x"e8",
          6410 => x"d6",
          6411 => x"ff",
          6412 => x"77",
          6413 => x"38",
          6414 => x"26",
          6415 => x"73",
          6416 => x"59",
          6417 => x"23",
          6418 => x"8b",
          6419 => x"ff",
          6420 => x"81",
          6421 => x"81",
          6422 => x"77",
          6423 => x"74",
          6424 => x"2a",
          6425 => x"51",
          6426 => x"80",
          6427 => x"73",
          6428 => x"92",
          6429 => x"1a",
          6430 => x"23",
          6431 => x"81",
          6432 => x"53",
          6433 => x"ff",
          6434 => x"9d",
          6435 => x"38",
          6436 => x"e8",
          6437 => x"d8",
          6438 => x"06",
          6439 => x"2e",
          6440 => x"0b",
          6441 => x"a0",
          6442 => x"78",
          6443 => x"3f",
          6444 => x"08",
          6445 => x"d8",
          6446 => x"98",
          6447 => x"84",
          6448 => x"80",
          6449 => x"0c",
          6450 => x"d8",
          6451 => x"0d",
          6452 => x"0d",
          6453 => x"40",
          6454 => x"78",
          6455 => x"3f",
          6456 => x"08",
          6457 => x"d8",
          6458 => x"38",
          6459 => x"5f",
          6460 => x"ac",
          6461 => x"19",
          6462 => x"51",
          6463 => x"82",
          6464 => x"58",
          6465 => x"08",
          6466 => x"9c",
          6467 => x"33",
          6468 => x"86",
          6469 => x"82",
          6470 => x"17",
          6471 => x"70",
          6472 => x"56",
          6473 => x"1a",
          6474 => x"e5",
          6475 => x"38",
          6476 => x"70",
          6477 => x"54",
          6478 => x"8e",
          6479 => x"b2",
          6480 => x"2e",
          6481 => x"81",
          6482 => x"19",
          6483 => x"2a",
          6484 => x"51",
          6485 => x"82",
          6486 => x"86",
          6487 => x"06",
          6488 => x"80",
          6489 => x"8d",
          6490 => x"81",
          6491 => x"90",
          6492 => x"1d",
          6493 => x"5e",
          6494 => x"09",
          6495 => x"b9",
          6496 => x"33",
          6497 => x"2e",
          6498 => x"81",
          6499 => x"1f",
          6500 => x"52",
          6501 => x"3f",
          6502 => x"08",
          6503 => x"06",
          6504 => x"95",
          6505 => x"70",
          6506 => x"29",
          6507 => x"56",
          6508 => x"5a",
          6509 => x"1b",
          6510 => x"51",
          6511 => x"82",
          6512 => x"83",
          6513 => x"56",
          6514 => x"b1",
          6515 => x"fe",
          6516 => x"38",
          6517 => x"df",
          6518 => x"d6",
          6519 => x"10",
          6520 => x"53",
          6521 => x"59",
          6522 => x"a1",
          6523 => x"d6",
          6524 => x"09",
          6525 => x"c1",
          6526 => x"8b",
          6527 => x"ff",
          6528 => x"81",
          6529 => x"81",
          6530 => x"7b",
          6531 => x"38",
          6532 => x"86",
          6533 => x"06",
          6534 => x"79",
          6535 => x"38",
          6536 => x"8b",
          6537 => x"1d",
          6538 => x"54",
          6539 => x"ff",
          6540 => x"ff",
          6541 => x"84",
          6542 => x"54",
          6543 => x"39",
          6544 => x"76",
          6545 => x"3f",
          6546 => x"08",
          6547 => x"54",
          6548 => x"bb",
          6549 => x"33",
          6550 => x"73",
          6551 => x"53",
          6552 => x"9c",
          6553 => x"e5",
          6554 => x"d6",
          6555 => x"2e",
          6556 => x"ff",
          6557 => x"ac",
          6558 => x"52",
          6559 => x"81",
          6560 => x"d8",
          6561 => x"d6",
          6562 => x"2e",
          6563 => x"77",
          6564 => x"0c",
          6565 => x"04",
          6566 => x"64",
          6567 => x"12",
          6568 => x"06",
          6569 => x"86",
          6570 => x"b5",
          6571 => x"1d",
          6572 => x"56",
          6573 => x"80",
          6574 => x"81",
          6575 => x"16",
          6576 => x"55",
          6577 => x"8c",
          6578 => x"70",
          6579 => x"70",
          6580 => x"e4",
          6581 => x"80",
          6582 => x"81",
          6583 => x"80",
          6584 => x"38",
          6585 => x"ab",
          6586 => x"5b",
          6587 => x"7b",
          6588 => x"53",
          6589 => x"51",
          6590 => x"85",
          6591 => x"c6",
          6592 => x"77",
          6593 => x"ff",
          6594 => x"55",
          6595 => x"b4",
          6596 => x"ff",
          6597 => x"19",
          6598 => x"57",
          6599 => x"76",
          6600 => x"81",
          6601 => x"2a",
          6602 => x"51",
          6603 => x"73",
          6604 => x"38",
          6605 => x"a1",
          6606 => x"17",
          6607 => x"25",
          6608 => x"39",
          6609 => x"02",
          6610 => x"05",
          6611 => x"b0",
          6612 => x"54",
          6613 => x"84",
          6614 => x"54",
          6615 => x"ff",
          6616 => x"76",
          6617 => x"58",
          6618 => x"38",
          6619 => x"05",
          6620 => x"fe",
          6621 => x"77",
          6622 => x"78",
          6623 => x"a0",
          6624 => x"74",
          6625 => x"52",
          6626 => x"3f",
          6627 => x"08",
          6628 => x"38",
          6629 => x"74",
          6630 => x"38",
          6631 => x"81",
          6632 => x"77",
          6633 => x"74",
          6634 => x"51",
          6635 => x"94",
          6636 => x"eb",
          6637 => x"15",
          6638 => x"58",
          6639 => x"87",
          6640 => x"81",
          6641 => x"70",
          6642 => x"57",
          6643 => x"87",
          6644 => x"38",
          6645 => x"f9",
          6646 => x"d8",
          6647 => x"81",
          6648 => x"e3",
          6649 => x"84",
          6650 => x"7a",
          6651 => x"82",
          6652 => x"d6",
          6653 => x"82",
          6654 => x"84",
          6655 => x"06",
          6656 => x"02",
          6657 => x"33",
          6658 => x"02",
          6659 => x"33",
          6660 => x"70",
          6661 => x"55",
          6662 => x"73",
          6663 => x"38",
          6664 => x"1d",
          6665 => x"86",
          6666 => x"d8",
          6667 => x"78",
          6668 => x"f3",
          6669 => x"d6",
          6670 => x"82",
          6671 => x"82",
          6672 => x"19",
          6673 => x"2e",
          6674 => x"78",
          6675 => x"1b",
          6676 => x"53",
          6677 => x"ef",
          6678 => x"d6",
          6679 => x"82",
          6680 => x"81",
          6681 => x"1a",
          6682 => x"3f",
          6683 => x"08",
          6684 => x"5d",
          6685 => x"52",
          6686 => x"ab",
          6687 => x"d8",
          6688 => x"d6",
          6689 => x"d7",
          6690 => x"08",
          6691 => x"7a",
          6692 => x"5a",
          6693 => x"8d",
          6694 => x"0b",
          6695 => x"82",
          6696 => x"8c",
          6697 => x"d6",
          6698 => x"9a",
          6699 => x"df",
          6700 => x"29",
          6701 => x"55",
          6702 => x"ff",
          6703 => x"38",
          6704 => x"70",
          6705 => x"57",
          6706 => x"52",
          6707 => x"17",
          6708 => x"51",
          6709 => x"73",
          6710 => x"ff",
          6711 => x"17",
          6712 => x"27",
          6713 => x"83",
          6714 => x"8b",
          6715 => x"1b",
          6716 => x"54",
          6717 => x"77",
          6718 => x"58",
          6719 => x"81",
          6720 => x"34",
          6721 => x"51",
          6722 => x"82",
          6723 => x"57",
          6724 => x"08",
          6725 => x"ff",
          6726 => x"fe",
          6727 => x"1a",
          6728 => x"51",
          6729 => x"82",
          6730 => x"57",
          6731 => x"08",
          6732 => x"53",
          6733 => x"08",
          6734 => x"08",
          6735 => x"3f",
          6736 => x"1a",
          6737 => x"08",
          6738 => x"3f",
          6739 => x"ab",
          6740 => x"06",
          6741 => x"8c",
          6742 => x"0b",
          6743 => x"76",
          6744 => x"d6",
          6745 => x"3d",
          6746 => x"3d",
          6747 => x"08",
          6748 => x"ac",
          6749 => x"59",
          6750 => x"ff",
          6751 => x"72",
          6752 => x"ed",
          6753 => x"d6",
          6754 => x"82",
          6755 => x"80",
          6756 => x"15",
          6757 => x"51",
          6758 => x"82",
          6759 => x"54",
          6760 => x"08",
          6761 => x"15",
          6762 => x"73",
          6763 => x"83",
          6764 => x"15",
          6765 => x"a2",
          6766 => x"d8",
          6767 => x"51",
          6768 => x"82",
          6769 => x"54",
          6770 => x"08",
          6771 => x"38",
          6772 => x"09",
          6773 => x"38",
          6774 => x"82",
          6775 => x"88",
          6776 => x"f4",
          6777 => x"60",
          6778 => x"59",
          6779 => x"96",
          6780 => x"1c",
          6781 => x"83",
          6782 => x"1c",
          6783 => x"81",
          6784 => x"70",
          6785 => x"05",
          6786 => x"57",
          6787 => x"57",
          6788 => x"81",
          6789 => x"10",
          6790 => x"81",
          6791 => x"53",
          6792 => x"80",
          6793 => x"70",
          6794 => x"06",
          6795 => x"8f",
          6796 => x"38",
          6797 => x"df",
          6798 => x"96",
          6799 => x"79",
          6800 => x"54",
          6801 => x"7a",
          6802 => x"07",
          6803 => x"98",
          6804 => x"d8",
          6805 => x"ff",
          6806 => x"ff",
          6807 => x"38",
          6808 => x"a5",
          6809 => x"2a",
          6810 => x"34",
          6811 => x"34",
          6812 => x"39",
          6813 => x"30",
          6814 => x"80",
          6815 => x"25",
          6816 => x"54",
          6817 => x"85",
          6818 => x"9a",
          6819 => x"34",
          6820 => x"17",
          6821 => x"8c",
          6822 => x"10",
          6823 => x"51",
          6824 => x"fe",
          6825 => x"30",
          6826 => x"70",
          6827 => x"59",
          6828 => x"17",
          6829 => x"80",
          6830 => x"34",
          6831 => x"1a",
          6832 => x"9c",
          6833 => x"70",
          6834 => x"5b",
          6835 => x"a0",
          6836 => x"74",
          6837 => x"81",
          6838 => x"81",
          6839 => x"89",
          6840 => x"70",
          6841 => x"25",
          6842 => x"76",
          6843 => x"38",
          6844 => x"8b",
          6845 => x"70",
          6846 => x"34",
          6847 => x"74",
          6848 => x"05",
          6849 => x"17",
          6850 => x"27",
          6851 => x"77",
          6852 => x"53",
          6853 => x"14",
          6854 => x"33",
          6855 => x"87",
          6856 => x"38",
          6857 => x"19",
          6858 => x"80",
          6859 => x"73",
          6860 => x"55",
          6861 => x"80",
          6862 => x"38",
          6863 => x"19",
          6864 => x"33",
          6865 => x"54",
          6866 => x"26",
          6867 => x"1c",
          6868 => x"33",
          6869 => x"79",
          6870 => x"72",
          6871 => x"85",
          6872 => x"2a",
          6873 => x"06",
          6874 => x"2e",
          6875 => x"15",
          6876 => x"ff",
          6877 => x"74",
          6878 => x"05",
          6879 => x"19",
          6880 => x"19",
          6881 => x"59",
          6882 => x"ff",
          6883 => x"17",
          6884 => x"80",
          6885 => x"34",
          6886 => x"8c",
          6887 => x"53",
          6888 => x"72",
          6889 => x"9c",
          6890 => x"8b",
          6891 => x"19",
          6892 => x"08",
          6893 => x"53",
          6894 => x"82",
          6895 => x"78",
          6896 => x"51",
          6897 => x"82",
          6898 => x"86",
          6899 => x"13",
          6900 => x"3f",
          6901 => x"08",
          6902 => x"8e",
          6903 => x"f0",
          6904 => x"70",
          6905 => x"80",
          6906 => x"51",
          6907 => x"af",
          6908 => x"81",
          6909 => x"dc",
          6910 => x"74",
          6911 => x"38",
          6912 => x"08",
          6913 => x"aa",
          6914 => x"44",
          6915 => x"33",
          6916 => x"73",
          6917 => x"81",
          6918 => x"81",
          6919 => x"dc",
          6920 => x"70",
          6921 => x"07",
          6922 => x"73",
          6923 => x"88",
          6924 => x"70",
          6925 => x"73",
          6926 => x"38",
          6927 => x"ab",
          6928 => x"52",
          6929 => x"ee",
          6930 => x"d8",
          6931 => x"e1",
          6932 => x"7d",
          6933 => x"08",
          6934 => x"59",
          6935 => x"05",
          6936 => x"3f",
          6937 => x"08",
          6938 => x"b1",
          6939 => x"ff",
          6940 => x"d8",
          6941 => x"38",
          6942 => x"82",
          6943 => x"90",
          6944 => x"73",
          6945 => x"19",
          6946 => x"d8",
          6947 => x"ff",
          6948 => x"32",
          6949 => x"73",
          6950 => x"25",
          6951 => x"55",
          6952 => x"38",
          6953 => x"2e",
          6954 => x"80",
          6955 => x"38",
          6956 => x"c6",
          6957 => x"92",
          6958 => x"d8",
          6959 => x"38",
          6960 => x"26",
          6961 => x"78",
          6962 => x"75",
          6963 => x"19",
          6964 => x"39",
          6965 => x"80",
          6966 => x"56",
          6967 => x"af",
          6968 => x"06",
          6969 => x"57",
          6970 => x"32",
          6971 => x"80",
          6972 => x"51",
          6973 => x"dc",
          6974 => x"9f",
          6975 => x"2b",
          6976 => x"2e",
          6977 => x"8c",
          6978 => x"54",
          6979 => x"a5",
          6980 => x"39",
          6981 => x"09",
          6982 => x"c9",
          6983 => x"22",
          6984 => x"2e",
          6985 => x"80",
          6986 => x"22",
          6987 => x"2e",
          6988 => x"b6",
          6989 => x"1a",
          6990 => x"23",
          6991 => x"1f",
          6992 => x"54",
          6993 => x"83",
          6994 => x"73",
          6995 => x"05",
          6996 => x"18",
          6997 => x"27",
          6998 => x"a0",
          6999 => x"ab",
          7000 => x"c4",
          7001 => x"2e",
          7002 => x"10",
          7003 => x"55",
          7004 => x"16",
          7005 => x"32",
          7006 => x"9f",
          7007 => x"53",
          7008 => x"75",
          7009 => x"38",
          7010 => x"ff",
          7011 => x"e0",
          7012 => x"7a",
          7013 => x"80",
          7014 => x"8d",
          7015 => x"85",
          7016 => x"83",
          7017 => x"99",
          7018 => x"22",
          7019 => x"ff",
          7020 => x"5d",
          7021 => x"09",
          7022 => x"38",
          7023 => x"10",
          7024 => x"51",
          7025 => x"a0",
          7026 => x"7c",
          7027 => x"83",
          7028 => x"54",
          7029 => x"09",
          7030 => x"38",
          7031 => x"57",
          7032 => x"aa",
          7033 => x"fe",
          7034 => x"51",
          7035 => x"2e",
          7036 => x"10",
          7037 => x"55",
          7038 => x"78",
          7039 => x"38",
          7040 => x"22",
          7041 => x"ae",
          7042 => x"06",
          7043 => x"53",
          7044 => x"1e",
          7045 => x"3f",
          7046 => x"5c",
          7047 => x"10",
          7048 => x"81",
          7049 => x"54",
          7050 => x"82",
          7051 => x"a0",
          7052 => x"75",
          7053 => x"30",
          7054 => x"51",
          7055 => x"79",
          7056 => x"73",
          7057 => x"38",
          7058 => x"57",
          7059 => x"54",
          7060 => x"78",
          7061 => x"81",
          7062 => x"32",
          7063 => x"72",
          7064 => x"70",
          7065 => x"51",
          7066 => x"80",
          7067 => x"7e",
          7068 => x"ae",
          7069 => x"2e",
          7070 => x"83",
          7071 => x"79",
          7072 => x"38",
          7073 => x"58",
          7074 => x"2b",
          7075 => x"5d",
          7076 => x"39",
          7077 => x"27",
          7078 => x"82",
          7079 => x"b5",
          7080 => x"80",
          7081 => x"82",
          7082 => x"83",
          7083 => x"70",
          7084 => x"81",
          7085 => x"56",
          7086 => x"8c",
          7087 => x"ff",
          7088 => x"e4",
          7089 => x"54",
          7090 => x"27",
          7091 => x"1f",
          7092 => x"26",
          7093 => x"83",
          7094 => x"57",
          7095 => x"7d",
          7096 => x"76",
          7097 => x"55",
          7098 => x"81",
          7099 => x"c3",
          7100 => x"2e",
          7101 => x"52",
          7102 => x"51",
          7103 => x"82",
          7104 => x"80",
          7105 => x"80",
          7106 => x"07",
          7107 => x"39",
          7108 => x"54",
          7109 => x"85",
          7110 => x"07",
          7111 => x"16",
          7112 => x"26",
          7113 => x"81",
          7114 => x"70",
          7115 => x"06",
          7116 => x"7d",
          7117 => x"54",
          7118 => x"81",
          7119 => x"de",
          7120 => x"33",
          7121 => x"e5",
          7122 => x"06",
          7123 => x"0b",
          7124 => x"7e",
          7125 => x"81",
          7126 => x"7b",
          7127 => x"fc",
          7128 => x"8c",
          7129 => x"8c",
          7130 => x"7b",
          7131 => x"73",
          7132 => x"81",
          7133 => x"76",
          7134 => x"76",
          7135 => x"81",
          7136 => x"73",
          7137 => x"81",
          7138 => x"80",
          7139 => x"76",
          7140 => x"7b",
          7141 => x"81",
          7142 => x"73",
          7143 => x"38",
          7144 => x"57",
          7145 => x"34",
          7146 => x"a5",
          7147 => x"d8",
          7148 => x"33",
          7149 => x"d6",
          7150 => x"2e",
          7151 => x"d6",
          7152 => x"2e",
          7153 => x"80",
          7154 => x"85",
          7155 => x"06",
          7156 => x"57",
          7157 => x"80",
          7158 => x"74",
          7159 => x"73",
          7160 => x"ed",
          7161 => x"0b",
          7162 => x"80",
          7163 => x"39",
          7164 => x"54",
          7165 => x"85",
          7166 => x"74",
          7167 => x"81",
          7168 => x"73",
          7169 => x"1e",
          7170 => x"2a",
          7171 => x"51",
          7172 => x"80",
          7173 => x"90",
          7174 => x"ff",
          7175 => x"b8",
          7176 => x"51",
          7177 => x"82",
          7178 => x"88",
          7179 => x"a1",
          7180 => x"d6",
          7181 => x"3d",
          7182 => x"3d",
          7183 => x"ff",
          7184 => x"71",
          7185 => x"5c",
          7186 => x"80",
          7187 => x"38",
          7188 => x"05",
          7189 => x"9f",
          7190 => x"71",
          7191 => x"38",
          7192 => x"71",
          7193 => x"81",
          7194 => x"38",
          7195 => x"11",
          7196 => x"06",
          7197 => x"70",
          7198 => x"38",
          7199 => x"81",
          7200 => x"05",
          7201 => x"76",
          7202 => x"38",
          7203 => x"c7",
          7204 => x"77",
          7205 => x"57",
          7206 => x"05",
          7207 => x"70",
          7208 => x"33",
          7209 => x"53",
          7210 => x"99",
          7211 => x"e0",
          7212 => x"ff",
          7213 => x"ff",
          7214 => x"70",
          7215 => x"38",
          7216 => x"81",
          7217 => x"51",
          7218 => x"9f",
          7219 => x"72",
          7220 => x"81",
          7221 => x"70",
          7222 => x"72",
          7223 => x"32",
          7224 => x"72",
          7225 => x"73",
          7226 => x"53",
          7227 => x"70",
          7228 => x"38",
          7229 => x"19",
          7230 => x"75",
          7231 => x"38",
          7232 => x"83",
          7233 => x"74",
          7234 => x"59",
          7235 => x"39",
          7236 => x"33",
          7237 => x"d6",
          7238 => x"3d",
          7239 => x"3d",
          7240 => x"80",
          7241 => x"34",
          7242 => x"17",
          7243 => x"75",
          7244 => x"3f",
          7245 => x"d6",
          7246 => x"80",
          7247 => x"16",
          7248 => x"3f",
          7249 => x"08",
          7250 => x"06",
          7251 => x"73",
          7252 => x"2e",
          7253 => x"80",
          7254 => x"0b",
          7255 => x"56",
          7256 => x"e9",
          7257 => x"06",
          7258 => x"57",
          7259 => x"32",
          7260 => x"80",
          7261 => x"51",
          7262 => x"8a",
          7263 => x"e8",
          7264 => x"06",
          7265 => x"53",
          7266 => x"52",
          7267 => x"51",
          7268 => x"82",
          7269 => x"55",
          7270 => x"08",
          7271 => x"38",
          7272 => x"c7",
          7273 => x"8a",
          7274 => x"ed",
          7275 => x"d8",
          7276 => x"d6",
          7277 => x"2e",
          7278 => x"55",
          7279 => x"d8",
          7280 => x"0d",
          7281 => x"0d",
          7282 => x"05",
          7283 => x"33",
          7284 => x"75",
          7285 => x"fc",
          7286 => x"d6",
          7287 => x"8b",
          7288 => x"82",
          7289 => x"24",
          7290 => x"82",
          7291 => x"84",
          7292 => x"a0",
          7293 => x"55",
          7294 => x"73",
          7295 => x"ee",
          7296 => x"0c",
          7297 => x"06",
          7298 => x"57",
          7299 => x"ae",
          7300 => x"33",
          7301 => x"3f",
          7302 => x"08",
          7303 => x"70",
          7304 => x"55",
          7305 => x"76",
          7306 => x"c0",
          7307 => x"2a",
          7308 => x"51",
          7309 => x"72",
          7310 => x"86",
          7311 => x"74",
          7312 => x"15",
          7313 => x"81",
          7314 => x"c6",
          7315 => x"d6",
          7316 => x"ff",
          7317 => x"06",
          7318 => x"56",
          7319 => x"38",
          7320 => x"8f",
          7321 => x"2a",
          7322 => x"51",
          7323 => x"72",
          7324 => x"80",
          7325 => x"52",
          7326 => x"3f",
          7327 => x"08",
          7328 => x"57",
          7329 => x"09",
          7330 => x"e2",
          7331 => x"74",
          7332 => x"56",
          7333 => x"33",
          7334 => x"72",
          7335 => x"38",
          7336 => x"51",
          7337 => x"82",
          7338 => x"57",
          7339 => x"84",
          7340 => x"ff",
          7341 => x"56",
          7342 => x"25",
          7343 => x"0b",
          7344 => x"56",
          7345 => x"05",
          7346 => x"83",
          7347 => x"2e",
          7348 => x"52",
          7349 => x"c6",
          7350 => x"d8",
          7351 => x"06",
          7352 => x"27",
          7353 => x"16",
          7354 => x"27",
          7355 => x"56",
          7356 => x"84",
          7357 => x"56",
          7358 => x"84",
          7359 => x"c3",
          7360 => x"c9",
          7361 => x"d8",
          7362 => x"ff",
          7363 => x"84",
          7364 => x"81",
          7365 => x"38",
          7366 => x"51",
          7367 => x"82",
          7368 => x"83",
          7369 => x"58",
          7370 => x"80",
          7371 => x"ca",
          7372 => x"d6",
          7373 => x"77",
          7374 => x"80",
          7375 => x"82",
          7376 => x"c8",
          7377 => x"11",
          7378 => x"06",
          7379 => x"8d",
          7380 => x"26",
          7381 => x"74",
          7382 => x"78",
          7383 => x"c5",
          7384 => x"59",
          7385 => x"15",
          7386 => x"2e",
          7387 => x"13",
          7388 => x"72",
          7389 => x"38",
          7390 => x"f2",
          7391 => x"14",
          7392 => x"3f",
          7393 => x"08",
          7394 => x"d8",
          7395 => x"23",
          7396 => x"57",
          7397 => x"83",
          7398 => x"cb",
          7399 => x"ad",
          7400 => x"d8",
          7401 => x"ff",
          7402 => x"8d",
          7403 => x"14",
          7404 => x"3f",
          7405 => x"08",
          7406 => x"14",
          7407 => x"3f",
          7408 => x"08",
          7409 => x"06",
          7410 => x"72",
          7411 => x"9e",
          7412 => x"22",
          7413 => x"84",
          7414 => x"5a",
          7415 => x"83",
          7416 => x"14",
          7417 => x"79",
          7418 => x"e0",
          7419 => x"d6",
          7420 => x"82",
          7421 => x"80",
          7422 => x"38",
          7423 => x"08",
          7424 => x"ff",
          7425 => x"38",
          7426 => x"83",
          7427 => x"83",
          7428 => x"74",
          7429 => x"85",
          7430 => x"89",
          7431 => x"76",
          7432 => x"ca",
          7433 => x"70",
          7434 => x"7b",
          7435 => x"73",
          7436 => x"17",
          7437 => x"b0",
          7438 => x"55",
          7439 => x"09",
          7440 => x"38",
          7441 => x"51",
          7442 => x"82",
          7443 => x"83",
          7444 => x"53",
          7445 => x"82",
          7446 => x"82",
          7447 => x"e4",
          7448 => x"80",
          7449 => x"d8",
          7450 => x"0c",
          7451 => x"53",
          7452 => x"56",
          7453 => x"81",
          7454 => x"13",
          7455 => x"74",
          7456 => x"82",
          7457 => x"74",
          7458 => x"81",
          7459 => x"06",
          7460 => x"83",
          7461 => x"2a",
          7462 => x"72",
          7463 => x"26",
          7464 => x"ff",
          7465 => x"0c",
          7466 => x"15",
          7467 => x"0b",
          7468 => x"76",
          7469 => x"81",
          7470 => x"38",
          7471 => x"51",
          7472 => x"82",
          7473 => x"83",
          7474 => x"53",
          7475 => x"09",
          7476 => x"f9",
          7477 => x"52",
          7478 => x"cb",
          7479 => x"d8",
          7480 => x"38",
          7481 => x"08",
          7482 => x"84",
          7483 => x"c6",
          7484 => x"d6",
          7485 => x"ff",
          7486 => x"72",
          7487 => x"2e",
          7488 => x"80",
          7489 => x"14",
          7490 => x"3f",
          7491 => x"08",
          7492 => x"a4",
          7493 => x"81",
          7494 => x"84",
          7495 => x"c6",
          7496 => x"d6",
          7497 => x"8a",
          7498 => x"2e",
          7499 => x"9d",
          7500 => x"14",
          7501 => x"3f",
          7502 => x"08",
          7503 => x"84",
          7504 => x"c6",
          7505 => x"d6",
          7506 => x"15",
          7507 => x"34",
          7508 => x"22",
          7509 => x"72",
          7510 => x"23",
          7511 => x"23",
          7512 => x"0b",
          7513 => x"80",
          7514 => x"0c",
          7515 => x"82",
          7516 => x"90",
          7517 => x"fb",
          7518 => x"54",
          7519 => x"80",
          7520 => x"73",
          7521 => x"80",
          7522 => x"72",
          7523 => x"80",
          7524 => x"86",
          7525 => x"15",
          7526 => x"71",
          7527 => x"81",
          7528 => x"81",
          7529 => x"ff",
          7530 => x"82",
          7531 => x"81",
          7532 => x"88",
          7533 => x"08",
          7534 => x"39",
          7535 => x"73",
          7536 => x"74",
          7537 => x"0c",
          7538 => x"04",
          7539 => x"02",
          7540 => x"7a",
          7541 => x"fc",
          7542 => x"f4",
          7543 => x"54",
          7544 => x"d6",
          7545 => x"bc",
          7546 => x"d8",
          7547 => x"82",
          7548 => x"70",
          7549 => x"73",
          7550 => x"38",
          7551 => x"78",
          7552 => x"2e",
          7553 => x"74",
          7554 => x"0c",
          7555 => x"80",
          7556 => x"80",
          7557 => x"70",
          7558 => x"51",
          7559 => x"82",
          7560 => x"54",
          7561 => x"d8",
          7562 => x"0d",
          7563 => x"0d",
          7564 => x"05",
          7565 => x"33",
          7566 => x"54",
          7567 => x"84",
          7568 => x"bf",
          7569 => x"99",
          7570 => x"53",
          7571 => x"05",
          7572 => x"f1",
          7573 => x"d8",
          7574 => x"d6",
          7575 => x"a4",
          7576 => x"69",
          7577 => x"70",
          7578 => x"f3",
          7579 => x"d8",
          7580 => x"d6",
          7581 => x"38",
          7582 => x"05",
          7583 => x"2b",
          7584 => x"80",
          7585 => x"86",
          7586 => x"06",
          7587 => x"2e",
          7588 => x"74",
          7589 => x"38",
          7590 => x"09",
          7591 => x"38",
          7592 => x"f4",
          7593 => x"d8",
          7594 => x"39",
          7595 => x"33",
          7596 => x"73",
          7597 => x"77",
          7598 => x"81",
          7599 => x"73",
          7600 => x"38",
          7601 => x"bc",
          7602 => x"07",
          7603 => x"b4",
          7604 => x"2a",
          7605 => x"51",
          7606 => x"2e",
          7607 => x"62",
          7608 => x"d7",
          7609 => x"d6",
          7610 => x"82",
          7611 => x"52",
          7612 => x"51",
          7613 => x"62",
          7614 => x"8b",
          7615 => x"53",
          7616 => x"51",
          7617 => x"80",
          7618 => x"05",
          7619 => x"3f",
          7620 => x"0b",
          7621 => x"75",
          7622 => x"f1",
          7623 => x"11",
          7624 => x"80",
          7625 => x"98",
          7626 => x"51",
          7627 => x"82",
          7628 => x"55",
          7629 => x"08",
          7630 => x"b7",
          7631 => x"c4",
          7632 => x"05",
          7633 => x"2a",
          7634 => x"51",
          7635 => x"80",
          7636 => x"84",
          7637 => x"39",
          7638 => x"70",
          7639 => x"54",
          7640 => x"a9",
          7641 => x"06",
          7642 => x"2e",
          7643 => x"55",
          7644 => x"73",
          7645 => x"c5",
          7646 => x"d6",
          7647 => x"ff",
          7648 => x"0c",
          7649 => x"d6",
          7650 => x"f8",
          7651 => x"2a",
          7652 => x"51",
          7653 => x"2e",
          7654 => x"80",
          7655 => x"7a",
          7656 => x"a0",
          7657 => x"a4",
          7658 => x"53",
          7659 => x"d5",
          7660 => x"d6",
          7661 => x"d6",
          7662 => x"1b",
          7663 => x"05",
          7664 => x"a0",
          7665 => x"d8",
          7666 => x"d8",
          7667 => x"0c",
          7668 => x"56",
          7669 => x"84",
          7670 => x"90",
          7671 => x"0b",
          7672 => x"80",
          7673 => x"0c",
          7674 => x"1a",
          7675 => x"2a",
          7676 => x"51",
          7677 => x"2e",
          7678 => x"82",
          7679 => x"80",
          7680 => x"38",
          7681 => x"08",
          7682 => x"8a",
          7683 => x"89",
          7684 => x"59",
          7685 => x"76",
          7686 => x"c6",
          7687 => x"d6",
          7688 => x"82",
          7689 => x"81",
          7690 => x"82",
          7691 => x"d8",
          7692 => x"09",
          7693 => x"38",
          7694 => x"78",
          7695 => x"30",
          7696 => x"80",
          7697 => x"77",
          7698 => x"38",
          7699 => x"06",
          7700 => x"c3",
          7701 => x"1a",
          7702 => x"38",
          7703 => x"06",
          7704 => x"2e",
          7705 => x"52",
          7706 => x"b1",
          7707 => x"d8",
          7708 => x"82",
          7709 => x"75",
          7710 => x"d6",
          7711 => x"9c",
          7712 => x"39",
          7713 => x"74",
          7714 => x"d6",
          7715 => x"3d",
          7716 => x"3d",
          7717 => x"65",
          7718 => x"5d",
          7719 => x"0c",
          7720 => x"05",
          7721 => x"f9",
          7722 => x"d6",
          7723 => x"82",
          7724 => x"8a",
          7725 => x"33",
          7726 => x"2e",
          7727 => x"56",
          7728 => x"90",
          7729 => x"06",
          7730 => x"74",
          7731 => x"b9",
          7732 => x"82",
          7733 => x"34",
          7734 => x"ad",
          7735 => x"91",
          7736 => x"56",
          7737 => x"8c",
          7738 => x"1a",
          7739 => x"74",
          7740 => x"38",
          7741 => x"80",
          7742 => x"38",
          7743 => x"70",
          7744 => x"56",
          7745 => x"b4",
          7746 => x"11",
          7747 => x"77",
          7748 => x"5b",
          7749 => x"38",
          7750 => x"88",
          7751 => x"8f",
          7752 => x"08",
          7753 => x"c4",
          7754 => x"d6",
          7755 => x"81",
          7756 => x"9f",
          7757 => x"2e",
          7758 => x"74",
          7759 => x"98",
          7760 => x"7e",
          7761 => x"3f",
          7762 => x"08",
          7763 => x"83",
          7764 => x"d8",
          7765 => x"89",
          7766 => x"77",
          7767 => x"d8",
          7768 => x"7f",
          7769 => x"58",
          7770 => x"75",
          7771 => x"75",
          7772 => x"77",
          7773 => x"7c",
          7774 => x"33",
          7775 => x"d4",
          7776 => x"d8",
          7777 => x"38",
          7778 => x"33",
          7779 => x"80",
          7780 => x"b4",
          7781 => x"31",
          7782 => x"27",
          7783 => x"80",
          7784 => x"52",
          7785 => x"77",
          7786 => x"7d",
          7787 => x"be",
          7788 => x"89",
          7789 => x"39",
          7790 => x"0c",
          7791 => x"83",
          7792 => x"80",
          7793 => x"55",
          7794 => x"83",
          7795 => x"9c",
          7796 => x"7e",
          7797 => x"3f",
          7798 => x"08",
          7799 => x"75",
          7800 => x"08",
          7801 => x"1f",
          7802 => x"7c",
          7803 => x"ec",
          7804 => x"31",
          7805 => x"7f",
          7806 => x"94",
          7807 => x"94",
          7808 => x"5c",
          7809 => x"80",
          7810 => x"d6",
          7811 => x"3d",
          7812 => x"3d",
          7813 => x"65",
          7814 => x"5d",
          7815 => x"0c",
          7816 => x"05",
          7817 => x"f6",
          7818 => x"d6",
          7819 => x"82",
          7820 => x"8a",
          7821 => x"33",
          7822 => x"2e",
          7823 => x"56",
          7824 => x"90",
          7825 => x"81",
          7826 => x"06",
          7827 => x"87",
          7828 => x"2e",
          7829 => x"95",
          7830 => x"91",
          7831 => x"56",
          7832 => x"81",
          7833 => x"34",
          7834 => x"94",
          7835 => x"08",
          7836 => x"56",
          7837 => x"84",
          7838 => x"5c",
          7839 => x"82",
          7840 => x"18",
          7841 => x"ff",
          7842 => x"74",
          7843 => x"7e",
          7844 => x"ff",
          7845 => x"2a",
          7846 => x"7a",
          7847 => x"8c",
          7848 => x"08",
          7849 => x"38",
          7850 => x"39",
          7851 => x"52",
          7852 => x"ef",
          7853 => x"d8",
          7854 => x"d6",
          7855 => x"2e",
          7856 => x"74",
          7857 => x"91",
          7858 => x"2e",
          7859 => x"74",
          7860 => x"88",
          7861 => x"38",
          7862 => x"0c",
          7863 => x"15",
          7864 => x"08",
          7865 => x"06",
          7866 => x"51",
          7867 => x"3f",
          7868 => x"08",
          7869 => x"98",
          7870 => x"7e",
          7871 => x"3f",
          7872 => x"08",
          7873 => x"d1",
          7874 => x"d8",
          7875 => x"89",
          7876 => x"78",
          7877 => x"d7",
          7878 => x"7f",
          7879 => x"58",
          7880 => x"75",
          7881 => x"75",
          7882 => x"78",
          7883 => x"7c",
          7884 => x"33",
          7885 => x"86",
          7886 => x"d8",
          7887 => x"38",
          7888 => x"08",
          7889 => x"56",
          7890 => x"9c",
          7891 => x"53",
          7892 => x"77",
          7893 => x"7d",
          7894 => x"16",
          7895 => x"fc",
          7896 => x"80",
          7897 => x"34",
          7898 => x"56",
          7899 => x"8c",
          7900 => x"19",
          7901 => x"38",
          7902 => x"bc",
          7903 => x"d6",
          7904 => x"df",
          7905 => x"b4",
          7906 => x"76",
          7907 => x"94",
          7908 => x"ff",
          7909 => x"71",
          7910 => x"7b",
          7911 => x"38",
          7912 => x"18",
          7913 => x"51",
          7914 => x"3f",
          7915 => x"08",
          7916 => x"75",
          7917 => x"94",
          7918 => x"ff",
          7919 => x"05",
          7920 => x"98",
          7921 => x"81",
          7922 => x"34",
          7923 => x"7e",
          7924 => x"0c",
          7925 => x"1a",
          7926 => x"94",
          7927 => x"1b",
          7928 => x"5e",
          7929 => x"27",
          7930 => x"55",
          7931 => x"0c",
          7932 => x"90",
          7933 => x"c0",
          7934 => x"90",
          7935 => x"56",
          7936 => x"d8",
          7937 => x"0d",
          7938 => x"0d",
          7939 => x"fc",
          7940 => x"52",
          7941 => x"3f",
          7942 => x"08",
          7943 => x"d8",
          7944 => x"38",
          7945 => x"70",
          7946 => x"81",
          7947 => x"55",
          7948 => x"80",
          7949 => x"16",
          7950 => x"51",
          7951 => x"3f",
          7952 => x"08",
          7953 => x"d8",
          7954 => x"38",
          7955 => x"8b",
          7956 => x"07",
          7957 => x"8b",
          7958 => x"16",
          7959 => x"52",
          7960 => x"cc",
          7961 => x"16",
          7962 => x"15",
          7963 => x"bd",
          7964 => x"b2",
          7965 => x"15",
          7966 => x"b1",
          7967 => x"92",
          7968 => x"b8",
          7969 => x"54",
          7970 => x"15",
          7971 => x"ff",
          7972 => x"82",
          7973 => x"90",
          7974 => x"bf",
          7975 => x"73",
          7976 => x"76",
          7977 => x"0c",
          7978 => x"04",
          7979 => x"76",
          7980 => x"fe",
          7981 => x"d6",
          7982 => x"82",
          7983 => x"9c",
          7984 => x"fc",
          7985 => x"51",
          7986 => x"82",
          7987 => x"53",
          7988 => x"08",
          7989 => x"d6",
          7990 => x"0c",
          7991 => x"d8",
          7992 => x"0d",
          7993 => x"0d",
          7994 => x"e6",
          7995 => x"52",
          7996 => x"d6",
          7997 => x"8b",
          7998 => x"d8",
          7999 => x"b4",
          8000 => x"71",
          8001 => x"0c",
          8002 => x"04",
          8003 => x"80",
          8004 => x"cc",
          8005 => x"3d",
          8006 => x"3f",
          8007 => x"08",
          8008 => x"d8",
          8009 => x"38",
          8010 => x"52",
          8011 => x"05",
          8012 => x"3f",
          8013 => x"08",
          8014 => x"d8",
          8015 => x"02",
          8016 => x"33",
          8017 => x"55",
          8018 => x"25",
          8019 => x"7a",
          8020 => x"54",
          8021 => x"a2",
          8022 => x"84",
          8023 => x"06",
          8024 => x"73",
          8025 => x"38",
          8026 => x"70",
          8027 => x"a5",
          8028 => x"d8",
          8029 => x"0c",
          8030 => x"d6",
          8031 => x"2e",
          8032 => x"83",
          8033 => x"74",
          8034 => x"0c",
          8035 => x"04",
          8036 => x"0d",
          8037 => x"08",
          8038 => x"08",
          8039 => x"7a",
          8040 => x"80",
          8041 => x"b4",
          8042 => x"e0",
          8043 => x"95",
          8044 => x"d8",
          8045 => x"d6",
          8046 => x"a1",
          8047 => x"d4",
          8048 => x"7c",
          8049 => x"80",
          8050 => x"55",
          8051 => x"3d",
          8052 => x"80",
          8053 => x"38",
          8054 => x"d3",
          8055 => x"55",
          8056 => x"82",
          8057 => x"57",
          8058 => x"08",
          8059 => x"80",
          8060 => x"52",
          8061 => x"b8",
          8062 => x"d6",
          8063 => x"82",
          8064 => x"82",
          8065 => x"da",
          8066 => x"7b",
          8067 => x"3f",
          8068 => x"08",
          8069 => x"0c",
          8070 => x"51",
          8071 => x"82",
          8072 => x"57",
          8073 => x"08",
          8074 => x"80",
          8075 => x"c9",
          8076 => x"d6",
          8077 => x"82",
          8078 => x"a7",
          8079 => x"3d",
          8080 => x"51",
          8081 => x"73",
          8082 => x"08",
          8083 => x"76",
          8084 => x"c5",
          8085 => x"d6",
          8086 => x"82",
          8087 => x"80",
          8088 => x"76",
          8089 => x"81",
          8090 => x"82",
          8091 => x"39",
          8092 => x"38",
          8093 => x"fd",
          8094 => x"74",
          8095 => x"3f",
          8096 => x"78",
          8097 => x"33",
          8098 => x"56",
          8099 => x"92",
          8100 => x"c6",
          8101 => x"16",
          8102 => x"33",
          8103 => x"73",
          8104 => x"16",
          8105 => x"26",
          8106 => x"75",
          8107 => x"38",
          8108 => x"05",
          8109 => x"80",
          8110 => x"11",
          8111 => x"18",
          8112 => x"58",
          8113 => x"34",
          8114 => x"ff",
          8115 => x"3d",
          8116 => x"58",
          8117 => x"fd",
          8118 => x"7b",
          8119 => x"06",
          8120 => x"18",
          8121 => x"08",
          8122 => x"af",
          8123 => x"0b",
          8124 => x"33",
          8125 => x"82",
          8126 => x"70",
          8127 => x"52",
          8128 => x"56",
          8129 => x"8d",
          8130 => x"70",
          8131 => x"51",
          8132 => x"f5",
          8133 => x"54",
          8134 => x"a7",
          8135 => x"74",
          8136 => x"38",
          8137 => x"73",
          8138 => x"81",
          8139 => x"81",
          8140 => x"39",
          8141 => x"81",
          8142 => x"74",
          8143 => x"81",
          8144 => x"91",
          8145 => x"80",
          8146 => x"18",
          8147 => x"54",
          8148 => x"70",
          8149 => x"34",
          8150 => x"eb",
          8151 => x"34",
          8152 => x"d8",
          8153 => x"3d",
          8154 => x"3d",
          8155 => x"8d",
          8156 => x"54",
          8157 => x"55",
          8158 => x"82",
          8159 => x"53",
          8160 => x"08",
          8161 => x"91",
          8162 => x"72",
          8163 => x"8c",
          8164 => x"73",
          8165 => x"38",
          8166 => x"70",
          8167 => x"81",
          8168 => x"57",
          8169 => x"73",
          8170 => x"08",
          8171 => x"94",
          8172 => x"75",
          8173 => x"9b",
          8174 => x"11",
          8175 => x"2b",
          8176 => x"73",
          8177 => x"38",
          8178 => x"16",
          8179 => x"de",
          8180 => x"d8",
          8181 => x"78",
          8182 => x"55",
          8183 => x"ce",
          8184 => x"d8",
          8185 => x"96",
          8186 => x"70",
          8187 => x"94",
          8188 => x"71",
          8189 => x"08",
          8190 => x"53",
          8191 => x"15",
          8192 => x"a7",
          8193 => x"74",
          8194 => x"97",
          8195 => x"d8",
          8196 => x"d6",
          8197 => x"2e",
          8198 => x"82",
          8199 => x"ff",
          8200 => x"38",
          8201 => x"08",
          8202 => x"73",
          8203 => x"73",
          8204 => x"9f",
          8205 => x"27",
          8206 => x"75",
          8207 => x"16",
          8208 => x"17",
          8209 => x"33",
          8210 => x"70",
          8211 => x"55",
          8212 => x"80",
          8213 => x"73",
          8214 => x"ff",
          8215 => x"82",
          8216 => x"54",
          8217 => x"08",
          8218 => x"d6",
          8219 => x"a8",
          8220 => x"74",
          8221 => x"cf",
          8222 => x"d8",
          8223 => x"ff",
          8224 => x"81",
          8225 => x"38",
          8226 => x"9c",
          8227 => x"a7",
          8228 => x"16",
          8229 => x"39",
          8230 => x"16",
          8231 => x"75",
          8232 => x"53",
          8233 => x"ab",
          8234 => x"79",
          8235 => x"ed",
          8236 => x"d8",
          8237 => x"82",
          8238 => x"34",
          8239 => x"c4",
          8240 => x"91",
          8241 => x"53",
          8242 => x"89",
          8243 => x"d8",
          8244 => x"94",
          8245 => x"8c",
          8246 => x"27",
          8247 => x"8c",
          8248 => x"15",
          8249 => x"07",
          8250 => x"16",
          8251 => x"ff",
          8252 => x"80",
          8253 => x"77",
          8254 => x"2e",
          8255 => x"9c",
          8256 => x"53",
          8257 => x"d8",
          8258 => x"0d",
          8259 => x"0d",
          8260 => x"54",
          8261 => x"81",
          8262 => x"53",
          8263 => x"05",
          8264 => x"84",
          8265 => x"9d",
          8266 => x"d8",
          8267 => x"d6",
          8268 => x"eb",
          8269 => x"0c",
          8270 => x"51",
          8271 => x"82",
          8272 => x"55",
          8273 => x"08",
          8274 => x"ab",
          8275 => x"98",
          8276 => x"80",
          8277 => x"38",
          8278 => x"70",
          8279 => x"81",
          8280 => x"57",
          8281 => x"ae",
          8282 => x"08",
          8283 => x"c2",
          8284 => x"d6",
          8285 => x"17",
          8286 => x"86",
          8287 => x"17",
          8288 => x"75",
          8289 => x"ae",
          8290 => x"d8",
          8291 => x"84",
          8292 => x"06",
          8293 => x"55",
          8294 => x"80",
          8295 => x"80",
          8296 => x"54",
          8297 => x"d8",
          8298 => x"0d",
          8299 => x"0d",
          8300 => x"fc",
          8301 => x"52",
          8302 => x"3f",
          8303 => x"08",
          8304 => x"d6",
          8305 => x"0c",
          8306 => x"04",
          8307 => x"77",
          8308 => x"fc",
          8309 => x"53",
          8310 => x"9b",
          8311 => x"d8",
          8312 => x"d6",
          8313 => x"e1",
          8314 => x"38",
          8315 => x"08",
          8316 => x"ff",
          8317 => x"82",
          8318 => x"53",
          8319 => x"82",
          8320 => x"52",
          8321 => x"a3",
          8322 => x"d8",
          8323 => x"d6",
          8324 => x"2e",
          8325 => x"85",
          8326 => x"87",
          8327 => x"d8",
          8328 => x"74",
          8329 => x"cf",
          8330 => x"52",
          8331 => x"bd",
          8332 => x"d6",
          8333 => x"32",
          8334 => x"72",
          8335 => x"70",
          8336 => x"08",
          8337 => x"54",
          8338 => x"d6",
          8339 => x"3d",
          8340 => x"3d",
          8341 => x"80",
          8342 => x"70",
          8343 => x"52",
          8344 => x"3f",
          8345 => x"08",
          8346 => x"d8",
          8347 => x"65",
          8348 => x"d2",
          8349 => x"d6",
          8350 => x"82",
          8351 => x"a0",
          8352 => x"cb",
          8353 => x"98",
          8354 => x"73",
          8355 => x"38",
          8356 => x"39",
          8357 => x"88",
          8358 => x"75",
          8359 => x"3f",
          8360 => x"d8",
          8361 => x"0d",
          8362 => x"0d",
          8363 => x"5c",
          8364 => x"3d",
          8365 => x"93",
          8366 => x"89",
          8367 => x"d8",
          8368 => x"d6",
          8369 => x"82",
          8370 => x"0c",
          8371 => x"11",
          8372 => x"94",
          8373 => x"56",
          8374 => x"74",
          8375 => x"75",
          8376 => x"e6",
          8377 => x"81",
          8378 => x"5b",
          8379 => x"82",
          8380 => x"75",
          8381 => x"73",
          8382 => x"81",
          8383 => x"38",
          8384 => x"57",
          8385 => x"3d",
          8386 => x"ff",
          8387 => x"82",
          8388 => x"ff",
          8389 => x"82",
          8390 => x"81",
          8391 => x"82",
          8392 => x"30",
          8393 => x"d8",
          8394 => x"25",
          8395 => x"19",
          8396 => x"5a",
          8397 => x"08",
          8398 => x"38",
          8399 => x"a8",
          8400 => x"d6",
          8401 => x"58",
          8402 => x"77",
          8403 => x"7d",
          8404 => x"ad",
          8405 => x"d6",
          8406 => x"82",
          8407 => x"80",
          8408 => x"70",
          8409 => x"ff",
          8410 => x"56",
          8411 => x"2e",
          8412 => x"9e",
          8413 => x"51",
          8414 => x"3f",
          8415 => x"08",
          8416 => x"06",
          8417 => x"80",
          8418 => x"19",
          8419 => x"54",
          8420 => x"14",
          8421 => x"cc",
          8422 => x"d8",
          8423 => x"06",
          8424 => x"80",
          8425 => x"19",
          8426 => x"54",
          8427 => x"06",
          8428 => x"79",
          8429 => x"78",
          8430 => x"79",
          8431 => x"84",
          8432 => x"07",
          8433 => x"84",
          8434 => x"82",
          8435 => x"92",
          8436 => x"f9",
          8437 => x"8a",
          8438 => x"53",
          8439 => x"e3",
          8440 => x"d6",
          8441 => x"82",
          8442 => x"81",
          8443 => x"17",
          8444 => x"81",
          8445 => x"17",
          8446 => x"2a",
          8447 => x"51",
          8448 => x"55",
          8449 => x"81",
          8450 => x"17",
          8451 => x"8c",
          8452 => x"81",
          8453 => x"9c",
          8454 => x"d8",
          8455 => x"17",
          8456 => x"51",
          8457 => x"3f",
          8458 => x"08",
          8459 => x"0c",
          8460 => x"39",
          8461 => x"52",
          8462 => x"ae",
          8463 => x"d6",
          8464 => x"2e",
          8465 => x"83",
          8466 => x"82",
          8467 => x"81",
          8468 => x"06",
          8469 => x"56",
          8470 => x"a1",
          8471 => x"82",
          8472 => x"9c",
          8473 => x"95",
          8474 => x"08",
          8475 => x"d8",
          8476 => x"51",
          8477 => x"3f",
          8478 => x"08",
          8479 => x"08",
          8480 => x"90",
          8481 => x"c0",
          8482 => x"90",
          8483 => x"80",
          8484 => x"75",
          8485 => x"75",
          8486 => x"d6",
          8487 => x"3d",
          8488 => x"3d",
          8489 => x"a2",
          8490 => x"05",
          8491 => x"51",
          8492 => x"82",
          8493 => x"55",
          8494 => x"08",
          8495 => x"78",
          8496 => x"08",
          8497 => x"70",
          8498 => x"93",
          8499 => x"d8",
          8500 => x"d6",
          8501 => x"df",
          8502 => x"ff",
          8503 => x"85",
          8504 => x"06",
          8505 => x"86",
          8506 => x"cb",
          8507 => x"2b",
          8508 => x"24",
          8509 => x"02",
          8510 => x"33",
          8511 => x"58",
          8512 => x"76",
          8513 => x"6c",
          8514 => x"ff",
          8515 => x"82",
          8516 => x"74",
          8517 => x"81",
          8518 => x"56",
          8519 => x"80",
          8520 => x"54",
          8521 => x"08",
          8522 => x"2e",
          8523 => x"73",
          8524 => x"d8",
          8525 => x"52",
          8526 => x"52",
          8527 => x"f6",
          8528 => x"d8",
          8529 => x"d6",
          8530 => x"eb",
          8531 => x"d8",
          8532 => x"51",
          8533 => x"3f",
          8534 => x"08",
          8535 => x"d8",
          8536 => x"87",
          8537 => x"39",
          8538 => x"08",
          8539 => x"38",
          8540 => x"08",
          8541 => x"77",
          8542 => x"3f",
          8543 => x"08",
          8544 => x"08",
          8545 => x"d6",
          8546 => x"80",
          8547 => x"55",
          8548 => x"95",
          8549 => x"2e",
          8550 => x"53",
          8551 => x"51",
          8552 => x"3f",
          8553 => x"08",
          8554 => x"38",
          8555 => x"a9",
          8556 => x"d6",
          8557 => x"74",
          8558 => x"0c",
          8559 => x"04",
          8560 => x"82",
          8561 => x"ff",
          8562 => x"9b",
          8563 => x"f5",
          8564 => x"d8",
          8565 => x"d6",
          8566 => x"b7",
          8567 => x"6a",
          8568 => x"70",
          8569 => x"f7",
          8570 => x"d8",
          8571 => x"d6",
          8572 => x"38",
          8573 => x"9b",
          8574 => x"d8",
          8575 => x"09",
          8576 => x"8f",
          8577 => x"df",
          8578 => x"85",
          8579 => x"51",
          8580 => x"74",
          8581 => x"78",
          8582 => x"8a",
          8583 => x"57",
          8584 => x"3f",
          8585 => x"08",
          8586 => x"82",
          8587 => x"83",
          8588 => x"82",
          8589 => x"81",
          8590 => x"06",
          8591 => x"54",
          8592 => x"08",
          8593 => x"81",
          8594 => x"81",
          8595 => x"39",
          8596 => x"38",
          8597 => x"08",
          8598 => x"ff",
          8599 => x"82",
          8600 => x"54",
          8601 => x"08",
          8602 => x"8b",
          8603 => x"b8",
          8604 => x"a5",
          8605 => x"54",
          8606 => x"15",
          8607 => x"90",
          8608 => x"15",
          8609 => x"b2",
          8610 => x"ce",
          8611 => x"a4",
          8612 => x"53",
          8613 => x"53",
          8614 => x"b2",
          8615 => x"78",
          8616 => x"80",
          8617 => x"ff",
          8618 => x"78",
          8619 => x"80",
          8620 => x"7f",
          8621 => x"d8",
          8622 => x"ff",
          8623 => x"78",
          8624 => x"83",
          8625 => x"51",
          8626 => x"3f",
          8627 => x"08",
          8628 => x"d8",
          8629 => x"82",
          8630 => x"52",
          8631 => x"51",
          8632 => x"3f",
          8633 => x"52",
          8634 => x"b7",
          8635 => x"54",
          8636 => x"15",
          8637 => x"81",
          8638 => x"34",
          8639 => x"a6",
          8640 => x"d6",
          8641 => x"8b",
          8642 => x"75",
          8643 => x"ff",
          8644 => x"73",
          8645 => x"0c",
          8646 => x"04",
          8647 => x"ab",
          8648 => x"51",
          8649 => x"82",
          8650 => x"fe",
          8651 => x"ab",
          8652 => x"91",
          8653 => x"d8",
          8654 => x"d6",
          8655 => x"d8",
          8656 => x"ab",
          8657 => x"9e",
          8658 => x"58",
          8659 => x"82",
          8660 => x"55",
          8661 => x"08",
          8662 => x"02",
          8663 => x"33",
          8664 => x"54",
          8665 => x"82",
          8666 => x"53",
          8667 => x"52",
          8668 => x"80",
          8669 => x"a2",
          8670 => x"53",
          8671 => x"3d",
          8672 => x"ff",
          8673 => x"ac",
          8674 => x"73",
          8675 => x"3f",
          8676 => x"08",
          8677 => x"d8",
          8678 => x"63",
          8679 => x"2e",
          8680 => x"88",
          8681 => x"3d",
          8682 => x"38",
          8683 => x"e8",
          8684 => x"d8",
          8685 => x"09",
          8686 => x"bb",
          8687 => x"ff",
          8688 => x"82",
          8689 => x"55",
          8690 => x"08",
          8691 => x"68",
          8692 => x"aa",
          8693 => x"05",
          8694 => x"51",
          8695 => x"3f",
          8696 => x"33",
          8697 => x"8b",
          8698 => x"84",
          8699 => x"06",
          8700 => x"73",
          8701 => x"a0",
          8702 => x"8b",
          8703 => x"54",
          8704 => x"15",
          8705 => x"33",
          8706 => x"70",
          8707 => x"55",
          8708 => x"2e",
          8709 => x"6f",
          8710 => x"e1",
          8711 => x"78",
          8712 => x"f1",
          8713 => x"d8",
          8714 => x"51",
          8715 => x"3f",
          8716 => x"d6",
          8717 => x"2e",
          8718 => x"82",
          8719 => x"52",
          8720 => x"a3",
          8721 => x"d6",
          8722 => x"80",
          8723 => x"58",
          8724 => x"d8",
          8725 => x"38",
          8726 => x"54",
          8727 => x"09",
          8728 => x"38",
          8729 => x"52",
          8730 => x"b4",
          8731 => x"54",
          8732 => x"15",
          8733 => x"82",
          8734 => x"9c",
          8735 => x"c1",
          8736 => x"d6",
          8737 => x"82",
          8738 => x"8c",
          8739 => x"ff",
          8740 => x"82",
          8741 => x"55",
          8742 => x"d8",
          8743 => x"0d",
          8744 => x"0d",
          8745 => x"05",
          8746 => x"05",
          8747 => x"33",
          8748 => x"53",
          8749 => x"05",
          8750 => x"51",
          8751 => x"82",
          8752 => x"55",
          8753 => x"08",
          8754 => x"78",
          8755 => x"96",
          8756 => x"51",
          8757 => x"82",
          8758 => x"55",
          8759 => x"08",
          8760 => x"80",
          8761 => x"81",
          8762 => x"86",
          8763 => x"38",
          8764 => x"61",
          8765 => x"12",
          8766 => x"7a",
          8767 => x"51",
          8768 => x"74",
          8769 => x"78",
          8770 => x"83",
          8771 => x"51",
          8772 => x"3f",
          8773 => x"08",
          8774 => x"d6",
          8775 => x"3d",
          8776 => x"3d",
          8777 => x"82",
          8778 => x"cc",
          8779 => x"3d",
          8780 => x"3f",
          8781 => x"08",
          8782 => x"d8",
          8783 => x"38",
          8784 => x"52",
          8785 => x"05",
          8786 => x"3f",
          8787 => x"08",
          8788 => x"d8",
          8789 => x"02",
          8790 => x"33",
          8791 => x"54",
          8792 => x"a6",
          8793 => x"22",
          8794 => x"71",
          8795 => x"53",
          8796 => x"51",
          8797 => x"3f",
          8798 => x"0b",
          8799 => x"76",
          8800 => x"ea",
          8801 => x"d8",
          8802 => x"82",
          8803 => x"94",
          8804 => x"e9",
          8805 => x"6c",
          8806 => x"53",
          8807 => x"05",
          8808 => x"51",
          8809 => x"82",
          8810 => x"82",
          8811 => x"30",
          8812 => x"d8",
          8813 => x"25",
          8814 => x"79",
          8815 => x"86",
          8816 => x"75",
          8817 => x"73",
          8818 => x"fa",
          8819 => x"80",
          8820 => x"8d",
          8821 => x"54",
          8822 => x"3f",
          8823 => x"08",
          8824 => x"d8",
          8825 => x"38",
          8826 => x"51",
          8827 => x"3f",
          8828 => x"08",
          8829 => x"d8",
          8830 => x"82",
          8831 => x"82",
          8832 => x"65",
          8833 => x"78",
          8834 => x"7b",
          8835 => x"55",
          8836 => x"34",
          8837 => x"8a",
          8838 => x"38",
          8839 => x"1a",
          8840 => x"34",
          8841 => x"9e",
          8842 => x"70",
          8843 => x"51",
          8844 => x"a0",
          8845 => x"8e",
          8846 => x"2e",
          8847 => x"86",
          8848 => x"34",
          8849 => x"30",
          8850 => x"80",
          8851 => x"7a",
          8852 => x"c1",
          8853 => x"2e",
          8854 => x"a4",
          8855 => x"51",
          8856 => x"3f",
          8857 => x"08",
          8858 => x"d8",
          8859 => x"7b",
          8860 => x"55",
          8861 => x"73",
          8862 => x"38",
          8863 => x"73",
          8864 => x"38",
          8865 => x"15",
          8866 => x"ff",
          8867 => x"82",
          8868 => x"7b",
          8869 => x"d6",
          8870 => x"3d",
          8871 => x"3d",
          8872 => x"9c",
          8873 => x"05",
          8874 => x"51",
          8875 => x"82",
          8876 => x"82",
          8877 => x"56",
          8878 => x"d8",
          8879 => x"38",
          8880 => x"52",
          8881 => x"52",
          8882 => x"b3",
          8883 => x"70",
          8884 => x"56",
          8885 => x"81",
          8886 => x"57",
          8887 => x"ff",
          8888 => x"82",
          8889 => x"83",
          8890 => x"80",
          8891 => x"d6",
          8892 => x"95",
          8893 => x"b5",
          8894 => x"d8",
          8895 => x"e8",
          8896 => x"d8",
          8897 => x"ff",
          8898 => x"80",
          8899 => x"74",
          8900 => x"e4",
          8901 => x"b2",
          8902 => x"d8",
          8903 => x"81",
          8904 => x"88",
          8905 => x"26",
          8906 => x"39",
          8907 => x"86",
          8908 => x"81",
          8909 => x"ff",
          8910 => x"38",
          8911 => x"54",
          8912 => x"81",
          8913 => x"81",
          8914 => x"77",
          8915 => x"59",
          8916 => x"6d",
          8917 => x"55",
          8918 => x"26",
          8919 => x"8a",
          8920 => x"86",
          8921 => x"e5",
          8922 => x"38",
          8923 => x"99",
          8924 => x"05",
          8925 => x"70",
          8926 => x"73",
          8927 => x"81",
          8928 => x"ff",
          8929 => x"ed",
          8930 => x"80",
          8931 => x"90",
          8932 => x"55",
          8933 => x"3f",
          8934 => x"08",
          8935 => x"d8",
          8936 => x"38",
          8937 => x"51",
          8938 => x"3f",
          8939 => x"08",
          8940 => x"d8",
          8941 => x"75",
          8942 => x"66",
          8943 => x"34",
          8944 => x"82",
          8945 => x"84",
          8946 => x"06",
          8947 => x"80",
          8948 => x"2e",
          8949 => x"81",
          8950 => x"ff",
          8951 => x"82",
          8952 => x"54",
          8953 => x"08",
          8954 => x"53",
          8955 => x"08",
          8956 => x"ff",
          8957 => x"66",
          8958 => x"8b",
          8959 => x"53",
          8960 => x"51",
          8961 => x"3f",
          8962 => x"0b",
          8963 => x"78",
          8964 => x"da",
          8965 => x"d8",
          8966 => x"55",
          8967 => x"d8",
          8968 => x"0d",
          8969 => x"0d",
          8970 => x"88",
          8971 => x"05",
          8972 => x"fc",
          8973 => x"54",
          8974 => x"d2",
          8975 => x"d6",
          8976 => x"82",
          8977 => x"82",
          8978 => x"1a",
          8979 => x"82",
          8980 => x"80",
          8981 => x"8c",
          8982 => x"78",
          8983 => x"1a",
          8984 => x"2a",
          8985 => x"51",
          8986 => x"90",
          8987 => x"82",
          8988 => x"58",
          8989 => x"81",
          8990 => x"39",
          8991 => x"22",
          8992 => x"70",
          8993 => x"56",
          8994 => x"af",
          8995 => x"14",
          8996 => x"30",
          8997 => x"9f",
          8998 => x"d8",
          8999 => x"19",
          9000 => x"5a",
          9001 => x"81",
          9002 => x"38",
          9003 => x"77",
          9004 => x"82",
          9005 => x"56",
          9006 => x"74",
          9007 => x"ff",
          9008 => x"81",
          9009 => x"55",
          9010 => x"75",
          9011 => x"82",
          9012 => x"d8",
          9013 => x"ff",
          9014 => x"d6",
          9015 => x"2e",
          9016 => x"82",
          9017 => x"8e",
          9018 => x"56",
          9019 => x"09",
          9020 => x"38",
          9021 => x"59",
          9022 => x"77",
          9023 => x"06",
          9024 => x"87",
          9025 => x"39",
          9026 => x"ba",
          9027 => x"55",
          9028 => x"2e",
          9029 => x"15",
          9030 => x"2e",
          9031 => x"83",
          9032 => x"75",
          9033 => x"7e",
          9034 => x"94",
          9035 => x"d8",
          9036 => x"d6",
          9037 => x"ce",
          9038 => x"16",
          9039 => x"56",
          9040 => x"38",
          9041 => x"19",
          9042 => x"90",
          9043 => x"7d",
          9044 => x"38",
          9045 => x"0c",
          9046 => x"0c",
          9047 => x"80",
          9048 => x"73",
          9049 => x"9c",
          9050 => x"05",
          9051 => x"57",
          9052 => x"26",
          9053 => x"7b",
          9054 => x"0c",
          9055 => x"81",
          9056 => x"84",
          9057 => x"54",
          9058 => x"d8",
          9059 => x"0d",
          9060 => x"0d",
          9061 => x"88",
          9062 => x"05",
          9063 => x"54",
          9064 => x"c5",
          9065 => x"56",
          9066 => x"d6",
          9067 => x"8b",
          9068 => x"d6",
          9069 => x"29",
          9070 => x"05",
          9071 => x"55",
          9072 => x"84",
          9073 => x"34",
          9074 => x"08",
          9075 => x"5f",
          9076 => x"51",
          9077 => x"3f",
          9078 => x"08",
          9079 => x"70",
          9080 => x"57",
          9081 => x"8b",
          9082 => x"82",
          9083 => x"06",
          9084 => x"56",
          9085 => x"38",
          9086 => x"05",
          9087 => x"7e",
          9088 => x"9e",
          9089 => x"d8",
          9090 => x"67",
          9091 => x"2e",
          9092 => x"82",
          9093 => x"8b",
          9094 => x"75",
          9095 => x"80",
          9096 => x"81",
          9097 => x"2e",
          9098 => x"80",
          9099 => x"38",
          9100 => x"0a",
          9101 => x"ff",
          9102 => x"55",
          9103 => x"86",
          9104 => x"8a",
          9105 => x"89",
          9106 => x"2a",
          9107 => x"77",
          9108 => x"59",
          9109 => x"81",
          9110 => x"70",
          9111 => x"07",
          9112 => x"56",
          9113 => x"38",
          9114 => x"05",
          9115 => x"7e",
          9116 => x"ae",
          9117 => x"82",
          9118 => x"8a",
          9119 => x"83",
          9120 => x"06",
          9121 => x"08",
          9122 => x"74",
          9123 => x"41",
          9124 => x"56",
          9125 => x"8a",
          9126 => x"61",
          9127 => x"55",
          9128 => x"27",
          9129 => x"93",
          9130 => x"80",
          9131 => x"38",
          9132 => x"70",
          9133 => x"43",
          9134 => x"95",
          9135 => x"06",
          9136 => x"2e",
          9137 => x"77",
          9138 => x"74",
          9139 => x"83",
          9140 => x"06",
          9141 => x"82",
          9142 => x"2e",
          9143 => x"78",
          9144 => x"2e",
          9145 => x"80",
          9146 => x"ae",
          9147 => x"2a",
          9148 => x"82",
          9149 => x"56",
          9150 => x"2e",
          9151 => x"77",
          9152 => x"82",
          9153 => x"79",
          9154 => x"70",
          9155 => x"5a",
          9156 => x"86",
          9157 => x"27",
          9158 => x"52",
          9159 => x"aa",
          9160 => x"d6",
          9161 => x"29",
          9162 => x"70",
          9163 => x"55",
          9164 => x"0b",
          9165 => x"08",
          9166 => x"05",
          9167 => x"ff",
          9168 => x"27",
          9169 => x"88",
          9170 => x"ae",
          9171 => x"2a",
          9172 => x"82",
          9173 => x"56",
          9174 => x"2e",
          9175 => x"77",
          9176 => x"82",
          9177 => x"79",
          9178 => x"70",
          9179 => x"5a",
          9180 => x"86",
          9181 => x"27",
          9182 => x"52",
          9183 => x"a9",
          9184 => x"d6",
          9185 => x"84",
          9186 => x"d6",
          9187 => x"f5",
          9188 => x"81",
          9189 => x"d8",
          9190 => x"d6",
          9191 => x"71",
          9192 => x"83",
          9193 => x"5e",
          9194 => x"89",
          9195 => x"5c",
          9196 => x"1c",
          9197 => x"05",
          9198 => x"ff",
          9199 => x"70",
          9200 => x"31",
          9201 => x"57",
          9202 => x"83",
          9203 => x"06",
          9204 => x"1c",
          9205 => x"5c",
          9206 => x"1d",
          9207 => x"29",
          9208 => x"31",
          9209 => x"55",
          9210 => x"87",
          9211 => x"7c",
          9212 => x"7a",
          9213 => x"31",
          9214 => x"a8",
          9215 => x"d6",
          9216 => x"7d",
          9217 => x"81",
          9218 => x"82",
          9219 => x"83",
          9220 => x"80",
          9221 => x"87",
          9222 => x"81",
          9223 => x"fd",
          9224 => x"f8",
          9225 => x"2e",
          9226 => x"80",
          9227 => x"ff",
          9228 => x"d6",
          9229 => x"a0",
          9230 => x"38",
          9231 => x"74",
          9232 => x"86",
          9233 => x"fd",
          9234 => x"81",
          9235 => x"80",
          9236 => x"83",
          9237 => x"39",
          9238 => x"08",
          9239 => x"92",
          9240 => x"b8",
          9241 => x"59",
          9242 => x"27",
          9243 => x"86",
          9244 => x"55",
          9245 => x"09",
          9246 => x"38",
          9247 => x"f5",
          9248 => x"38",
          9249 => x"55",
          9250 => x"86",
          9251 => x"80",
          9252 => x"7a",
          9253 => x"e7",
          9254 => x"82",
          9255 => x"7a",
          9256 => x"b8",
          9257 => x"52",
          9258 => x"ff",
          9259 => x"79",
          9260 => x"7b",
          9261 => x"06",
          9262 => x"51",
          9263 => x"3f",
          9264 => x"1c",
          9265 => x"32",
          9266 => x"96",
          9267 => x"06",
          9268 => x"91",
          9269 => x"8f",
          9270 => x"55",
          9271 => x"ff",
          9272 => x"74",
          9273 => x"06",
          9274 => x"51",
          9275 => x"3f",
          9276 => x"52",
          9277 => x"ff",
          9278 => x"f8",
          9279 => x"34",
          9280 => x"1b",
          9281 => x"87",
          9282 => x"52",
          9283 => x"ff",
          9284 => x"60",
          9285 => x"51",
          9286 => x"3f",
          9287 => x"09",
          9288 => x"cb",
          9289 => x"b2",
          9290 => x"c3",
          9291 => x"8e",
          9292 => x"52",
          9293 => x"ff",
          9294 => x"82",
          9295 => x"51",
          9296 => x"3f",
          9297 => x"1b",
          9298 => x"c3",
          9299 => x"b2",
          9300 => x"8e",
          9301 => x"80",
          9302 => x"1c",
          9303 => x"80",
          9304 => x"93",
          9305 => x"9c",
          9306 => x"1b",
          9307 => x"82",
          9308 => x"52",
          9309 => x"ff",
          9310 => x"7c",
          9311 => x"06",
          9312 => x"51",
          9313 => x"3f",
          9314 => x"a4",
          9315 => x"0b",
          9316 => x"93",
          9317 => x"b0",
          9318 => x"51",
          9319 => x"3f",
          9320 => x"52",
          9321 => x"70",
          9322 => x"8d",
          9323 => x"54",
          9324 => x"52",
          9325 => x"8a",
          9326 => x"56",
          9327 => x"08",
          9328 => x"7d",
          9329 => x"81",
          9330 => x"38",
          9331 => x"86",
          9332 => x"52",
          9333 => x"89",
          9334 => x"80",
          9335 => x"7a",
          9336 => x"9b",
          9337 => x"85",
          9338 => x"7a",
          9339 => x"bd",
          9340 => x"85",
          9341 => x"83",
          9342 => x"ff",
          9343 => x"ff",
          9344 => x"e8",
          9345 => x"8d",
          9346 => x"52",
          9347 => x"51",
          9348 => x"3f",
          9349 => x"52",
          9350 => x"8c",
          9351 => x"54",
          9352 => x"53",
          9353 => x"51",
          9354 => x"3f",
          9355 => x"16",
          9356 => x"7e",
          9357 => x"86",
          9358 => x"80",
          9359 => x"ff",
          9360 => x"7f",
          9361 => x"7d",
          9362 => x"81",
          9363 => x"f8",
          9364 => x"ff",
          9365 => x"ff",
          9366 => x"51",
          9367 => x"3f",
          9368 => x"88",
          9369 => x"39",
          9370 => x"f8",
          9371 => x"2e",
          9372 => x"55",
          9373 => x"51",
          9374 => x"3f",
          9375 => x"57",
          9376 => x"83",
          9377 => x"76",
          9378 => x"7a",
          9379 => x"ff",
          9380 => x"82",
          9381 => x"82",
          9382 => x"80",
          9383 => x"d8",
          9384 => x"51",
          9385 => x"3f",
          9386 => x"78",
          9387 => x"74",
          9388 => x"18",
          9389 => x"2e",
          9390 => x"79",
          9391 => x"2e",
          9392 => x"55",
          9393 => x"62",
          9394 => x"74",
          9395 => x"75",
          9396 => x"7e",
          9397 => x"e6",
          9398 => x"d8",
          9399 => x"38",
          9400 => x"78",
          9401 => x"74",
          9402 => x"56",
          9403 => x"93",
          9404 => x"66",
          9405 => x"26",
          9406 => x"56",
          9407 => x"83",
          9408 => x"64",
          9409 => x"77",
          9410 => x"84",
          9411 => x"52",
          9412 => x"8b",
          9413 => x"d4",
          9414 => x"51",
          9415 => x"3f",
          9416 => x"55",
          9417 => x"81",
          9418 => x"34",
          9419 => x"16",
          9420 => x"16",
          9421 => x"16",
          9422 => x"05",
          9423 => x"c1",
          9424 => x"fe",
          9425 => x"fe",
          9426 => x"34",
          9427 => x"08",
          9428 => x"07",
          9429 => x"16",
          9430 => x"d8",
          9431 => x"34",
          9432 => x"c6",
          9433 => x"8a",
          9434 => x"52",
          9435 => x"51",
          9436 => x"3f",
          9437 => x"53",
          9438 => x"51",
          9439 => x"3f",
          9440 => x"d6",
          9441 => x"38",
          9442 => x"52",
          9443 => x"88",
          9444 => x"56",
          9445 => x"08",
          9446 => x"39",
          9447 => x"39",
          9448 => x"39",
          9449 => x"08",
          9450 => x"d6",
          9451 => x"3d",
          9452 => x"3d",
          9453 => x"5b",
          9454 => x"60",
          9455 => x"57",
          9456 => x"25",
          9457 => x"3d",
          9458 => x"55",
          9459 => x"15",
          9460 => x"c9",
          9461 => x"81",
          9462 => x"06",
          9463 => x"3d",
          9464 => x"8d",
          9465 => x"74",
          9466 => x"05",
          9467 => x"17",
          9468 => x"2e",
          9469 => x"c9",
          9470 => x"34",
          9471 => x"83",
          9472 => x"74",
          9473 => x"0c",
          9474 => x"04",
          9475 => x"7b",
          9476 => x"b3",
          9477 => x"57",
          9478 => x"09",
          9479 => x"38",
          9480 => x"51",
          9481 => x"17",
          9482 => x"76",
          9483 => x"88",
          9484 => x"17",
          9485 => x"59",
          9486 => x"81",
          9487 => x"76",
          9488 => x"8b",
          9489 => x"54",
          9490 => x"17",
          9491 => x"51",
          9492 => x"79",
          9493 => x"30",
          9494 => x"9f",
          9495 => x"53",
          9496 => x"75",
          9497 => x"81",
          9498 => x"0c",
          9499 => x"04",
          9500 => x"79",
          9501 => x"56",
          9502 => x"24",
          9503 => x"3d",
          9504 => x"74",
          9505 => x"52",
          9506 => x"cb",
          9507 => x"d6",
          9508 => x"38",
          9509 => x"78",
          9510 => x"06",
          9511 => x"16",
          9512 => x"39",
          9513 => x"82",
          9514 => x"89",
          9515 => x"fd",
          9516 => x"54",
          9517 => x"80",
          9518 => x"ff",
          9519 => x"76",
          9520 => x"3d",
          9521 => x"3d",
          9522 => x"e3",
          9523 => x"53",
          9524 => x"53",
          9525 => x"3f",
          9526 => x"51",
          9527 => x"72",
          9528 => x"3f",
          9529 => x"04",
          9530 => x"75",
          9531 => x"9a",
          9532 => x"53",
          9533 => x"80",
          9534 => x"38",
          9535 => x"ff",
          9536 => x"c3",
          9537 => x"ff",
          9538 => x"73",
          9539 => x"09",
          9540 => x"38",
          9541 => x"af",
          9542 => x"98",
          9543 => x"71",
          9544 => x"81",
          9545 => x"ff",
          9546 => x"51",
          9547 => x"26",
          9548 => x"10",
          9549 => x"05",
          9550 => x"51",
          9551 => x"80",
          9552 => x"ff",
          9553 => x"71",
          9554 => x"0c",
          9555 => x"04",
          9556 => x"02",
          9557 => x"02",
          9558 => x"05",
          9559 => x"80",
          9560 => x"ff",
          9561 => x"70",
          9562 => x"71",
          9563 => x"09",
          9564 => x"38",
          9565 => x"26",
          9566 => x"10",
          9567 => x"05",
          9568 => x"51",
          9569 => x"d8",
          9570 => x"0d",
          9571 => x"0d",
          9572 => x"83",
          9573 => x"81",
          9574 => x"83",
          9575 => x"82",
          9576 => x"52",
          9577 => x"27",
          9578 => x"cf",
          9579 => x"70",
          9580 => x"22",
          9581 => x"80",
          9582 => x"26",
          9583 => x"55",
          9584 => x"38",
          9585 => x"05",
          9586 => x"88",
          9587 => x"ff",
          9588 => x"54",
          9589 => x"71",
          9590 => x"d7",
          9591 => x"26",
          9592 => x"73",
          9593 => x"ae",
          9594 => x"70",
          9595 => x"75",
          9596 => x"11",
          9597 => x"51",
          9598 => x"39",
          9599 => x"81",
          9600 => x"31",
          9601 => x"39",
          9602 => x"9f",
          9603 => x"51",
          9604 => x"12",
          9605 => x"e6",
          9606 => x"39",
          9607 => x"8b",
          9608 => x"12",
          9609 => x"c7",
          9610 => x"70",
          9611 => x"06",
          9612 => x"73",
          9613 => x"72",
          9614 => x"fe",
          9615 => x"51",
          9616 => x"d8",
          9617 => x"0d",
          9618 => x"00",
          9619 => x"ff",
          9620 => x"ff",
          9621 => x"ff",
          9622 => x"00",
          9623 => x"51",
          9624 => x"d5",
          9625 => x"dc",
          9626 => x"e3",
          9627 => x"ea",
          9628 => x"f1",
          9629 => x"f8",
          9630 => x"ff",
          9631 => x"06",
          9632 => x"0d",
          9633 => x"14",
          9634 => x"1b",
          9635 => x"21",
          9636 => x"27",
          9637 => x"2d",
          9638 => x"33",
          9639 => x"39",
          9640 => x"3f",
          9641 => x"45",
          9642 => x"4b",
          9643 => x"34",
          9644 => x"3a",
          9645 => x"40",
          9646 => x"46",
          9647 => x"4c",
          9648 => x"2a",
          9649 => x"2a",
          9650 => x"3b",
          9651 => x"93",
          9652 => x"12",
          9653 => x"ff",
          9654 => x"03",
          9655 => x"64",
          9656 => x"46",
          9657 => x"dc",
          9658 => x"62",
          9659 => x"e5",
          9660 => x"ff",
          9661 => x"3b",
          9662 => x"64",
          9663 => x"03",
          9664 => x"ff",
          9665 => x"ff",
          9666 => x"62",
          9667 => x"dc",
          9668 => x"64",
          9669 => x"93",
          9670 => x"ee",
          9671 => x"fc",
          9672 => x"08",
          9673 => x"0d",
          9674 => x"12",
          9675 => x"17",
          9676 => x"1c",
          9677 => x"21",
          9678 => x"27",
          9679 => x"31",
          9680 => x"1a",
          9681 => x"1a",
          9682 => x"60",
          9683 => x"1a",
          9684 => x"1a",
          9685 => x"1a",
          9686 => x"1a",
          9687 => x"1a",
          9688 => x"1a",
          9689 => x"1a",
          9690 => x"1d",
          9691 => x"1a",
          9692 => x"48",
          9693 => x"78",
          9694 => x"1a",
          9695 => x"1a",
          9696 => x"1a",
          9697 => x"1a",
          9698 => x"1a",
          9699 => x"1a",
          9700 => x"1a",
          9701 => x"1a",
          9702 => x"1a",
          9703 => x"1a",
          9704 => x"1a",
          9705 => x"1a",
          9706 => x"1a",
          9707 => x"1a",
          9708 => x"1a",
          9709 => x"1a",
          9710 => x"1a",
          9711 => x"1a",
          9712 => x"1a",
          9713 => x"1a",
          9714 => x"1a",
          9715 => x"1a",
          9716 => x"1a",
          9717 => x"1a",
          9718 => x"1a",
          9719 => x"1a",
          9720 => x"1a",
          9721 => x"1a",
          9722 => x"1a",
          9723 => x"1a",
          9724 => x"1a",
          9725 => x"1a",
          9726 => x"1a",
          9727 => x"1a",
          9728 => x"1a",
          9729 => x"1a",
          9730 => x"a8",
          9731 => x"1a",
          9732 => x"1a",
          9733 => x"1a",
          9734 => x"1a",
          9735 => x"16",
          9736 => x"1a",
          9737 => x"1a",
          9738 => x"1a",
          9739 => x"1a",
          9740 => x"1a",
          9741 => x"1a",
          9742 => x"1a",
          9743 => x"1a",
          9744 => x"1a",
          9745 => x"1a",
          9746 => x"d8",
          9747 => x"3f",
          9748 => x"af",
          9749 => x"af",
          9750 => x"af",
          9751 => x"1a",
          9752 => x"3f",
          9753 => x"1a",
          9754 => x"1a",
          9755 => x"98",
          9756 => x"1a",
          9757 => x"1a",
          9758 => x"ec",
          9759 => x"f7",
          9760 => x"1a",
          9761 => x"1a",
          9762 => x"11",
          9763 => x"1a",
          9764 => x"1f",
          9765 => x"1a",
          9766 => x"1a",
          9767 => x"16",
          9768 => x"69",
          9769 => x"00",
          9770 => x"63",
          9771 => x"00",
          9772 => x"69",
          9773 => x"00",
          9774 => x"61",
          9775 => x"00",
          9776 => x"65",
          9777 => x"00",
          9778 => x"65",
          9779 => x"00",
          9780 => x"70",
          9781 => x"00",
          9782 => x"66",
          9783 => x"00",
          9784 => x"6d",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"6c",
          9794 => x"00",
          9795 => x"00",
          9796 => x"74",
          9797 => x"00",
          9798 => x"65",
          9799 => x"00",
          9800 => x"6f",
          9801 => x"00",
          9802 => x"74",
          9803 => x"00",
          9804 => x"73",
          9805 => x"00",
          9806 => x"73",
          9807 => x"00",
          9808 => x"6f",
          9809 => x"00",
          9810 => x"00",
          9811 => x"6b",
          9812 => x"72",
          9813 => x"00",
          9814 => x"65",
          9815 => x"6c",
          9816 => x"72",
          9817 => x"00",
          9818 => x"6b",
          9819 => x"74",
          9820 => x"61",
          9821 => x"00",
          9822 => x"66",
          9823 => x"20",
          9824 => x"6e",
          9825 => x"00",
          9826 => x"70",
          9827 => x"20",
          9828 => x"6e",
          9829 => x"00",
          9830 => x"61",
          9831 => x"20",
          9832 => x"65",
          9833 => x"65",
          9834 => x"00",
          9835 => x"65",
          9836 => x"64",
          9837 => x"65",
          9838 => x"00",
          9839 => x"65",
          9840 => x"72",
          9841 => x"79",
          9842 => x"69",
          9843 => x"2e",
          9844 => x"00",
          9845 => x"65",
          9846 => x"6e",
          9847 => x"20",
          9848 => x"61",
          9849 => x"2e",
          9850 => x"00",
          9851 => x"69",
          9852 => x"72",
          9853 => x"20",
          9854 => x"74",
          9855 => x"65",
          9856 => x"00",
          9857 => x"76",
          9858 => x"75",
          9859 => x"72",
          9860 => x"20",
          9861 => x"61",
          9862 => x"2e",
          9863 => x"00",
          9864 => x"6b",
          9865 => x"74",
          9866 => x"61",
          9867 => x"64",
          9868 => x"00",
          9869 => x"63",
          9870 => x"61",
          9871 => x"6c",
          9872 => x"69",
          9873 => x"79",
          9874 => x"6d",
          9875 => x"75",
          9876 => x"6f",
          9877 => x"69",
          9878 => x"00",
          9879 => x"6d",
          9880 => x"61",
          9881 => x"74",
          9882 => x"00",
          9883 => x"65",
          9884 => x"2c",
          9885 => x"65",
          9886 => x"69",
          9887 => x"63",
          9888 => x"65",
          9889 => x"64",
          9890 => x"00",
          9891 => x"65",
          9892 => x"20",
          9893 => x"6b",
          9894 => x"00",
          9895 => x"75",
          9896 => x"63",
          9897 => x"74",
          9898 => x"6d",
          9899 => x"2e",
          9900 => x"00",
          9901 => x"20",
          9902 => x"79",
          9903 => x"65",
          9904 => x"69",
          9905 => x"2e",
          9906 => x"00",
          9907 => x"61",
          9908 => x"65",
          9909 => x"69",
          9910 => x"72",
          9911 => x"74",
          9912 => x"00",
          9913 => x"63",
          9914 => x"2e",
          9915 => x"00",
          9916 => x"6e",
          9917 => x"20",
          9918 => x"6f",
          9919 => x"00",
          9920 => x"75",
          9921 => x"74",
          9922 => x"25",
          9923 => x"74",
          9924 => x"75",
          9925 => x"74",
          9926 => x"73",
          9927 => x"0a",
          9928 => x"00",
          9929 => x"64",
          9930 => x"00",
          9931 => x"30",
          9932 => x"2c",
          9933 => x"25",
          9934 => x"78",
          9935 => x"3d",
          9936 => x"6c",
          9937 => x"5f",
          9938 => x"3d",
          9939 => x"6c",
          9940 => x"30",
          9941 => x"20",
          9942 => x"6c",
          9943 => x"00",
          9944 => x"6c",
          9945 => x"00",
          9946 => x"00",
          9947 => x"58",
          9948 => x"00",
          9949 => x"20",
          9950 => x"20",
          9951 => x"00",
          9952 => x"58",
          9953 => x"00",
          9954 => x"00",
          9955 => x"00",
          9956 => x"00",
          9957 => x"00",
          9958 => x"20",
          9959 => x"28",
          9960 => x"00",
          9961 => x"31",
          9962 => x"30",
          9963 => x"00",
          9964 => x"30",
          9965 => x"00",
          9966 => x"55",
          9967 => x"65",
          9968 => x"30",
          9969 => x"20",
          9970 => x"25",
          9971 => x"2a",
          9972 => x"00",
          9973 => x"20",
          9974 => x"65",
          9975 => x"70",
          9976 => x"61",
          9977 => x"65",
          9978 => x"00",
          9979 => x"65",
          9980 => x"6e",
          9981 => x"72",
          9982 => x"00",
          9983 => x"20",
          9984 => x"65",
          9985 => x"70",
          9986 => x"00",
          9987 => x"54",
          9988 => x"44",
          9989 => x"74",
          9990 => x"75",
          9991 => x"00",
          9992 => x"54",
          9993 => x"52",
          9994 => x"74",
          9995 => x"75",
          9996 => x"00",
          9997 => x"54",
          9998 => x"58",
          9999 => x"74",
         10000 => x"75",
         10001 => x"00",
         10002 => x"54",
         10003 => x"58",
         10004 => x"74",
         10005 => x"75",
         10006 => x"00",
         10007 => x"54",
         10008 => x"58",
         10009 => x"74",
         10010 => x"75",
         10011 => x"00",
         10012 => x"54",
         10013 => x"58",
         10014 => x"74",
         10015 => x"75",
         10016 => x"00",
         10017 => x"74",
         10018 => x"20",
         10019 => x"74",
         10020 => x"72",
         10021 => x"00",
         10022 => x"62",
         10023 => x"67",
         10024 => x"6d",
         10025 => x"2e",
         10026 => x"00",
         10027 => x"6f",
         10028 => x"63",
         10029 => x"74",
         10030 => x"00",
         10031 => x"2e",
         10032 => x"00",
         10033 => x"00",
         10034 => x"6c",
         10035 => x"74",
         10036 => x"6e",
         10037 => x"61",
         10038 => x"65",
         10039 => x"20",
         10040 => x"64",
         10041 => x"20",
         10042 => x"61",
         10043 => x"69",
         10044 => x"20",
         10045 => x"75",
         10046 => x"79",
         10047 => x"00",
         10048 => x"00",
         10049 => x"61",
         10050 => x"67",
         10051 => x"2e",
         10052 => x"00",
         10053 => x"79",
         10054 => x"2e",
         10055 => x"00",
         10056 => x"70",
         10057 => x"6e",
         10058 => x"2e",
         10059 => x"00",
         10060 => x"6c",
         10061 => x"30",
         10062 => x"2d",
         10063 => x"38",
         10064 => x"25",
         10065 => x"29",
         10066 => x"00",
         10067 => x"70",
         10068 => x"6d",
         10069 => x"00",
         10070 => x"6d",
         10071 => x"74",
         10072 => x"00",
         10073 => x"6c",
         10074 => x"30",
         10075 => x"00",
         10076 => x"00",
         10077 => x"6c",
         10078 => x"30",
         10079 => x"00",
         10080 => x"6c",
         10081 => x"30",
         10082 => x"2d",
         10083 => x"00",
         10084 => x"63",
         10085 => x"6e",
         10086 => x"6f",
         10087 => x"40",
         10088 => x"38",
         10089 => x"2e",
         10090 => x"00",
         10091 => x"6c",
         10092 => x"20",
         10093 => x"65",
         10094 => x"25",
         10095 => x"78",
         10096 => x"2e",
         10097 => x"00",
         10098 => x"6c",
         10099 => x"74",
         10100 => x"65",
         10101 => x"6f",
         10102 => x"28",
         10103 => x"2e",
         10104 => x"00",
         10105 => x"74",
         10106 => x"69",
         10107 => x"61",
         10108 => x"69",
         10109 => x"69",
         10110 => x"2e",
         10111 => x"00",
         10112 => x"64",
         10113 => x"62",
         10114 => x"69",
         10115 => x"2e",
         10116 => x"00",
         10117 => x"00",
         10118 => x"00",
         10119 => x"5c",
         10120 => x"25",
         10121 => x"73",
         10122 => x"00",
         10123 => x"5c",
         10124 => x"25",
         10125 => x"00",
         10126 => x"5c",
         10127 => x"00",
         10128 => x"20",
         10129 => x"6d",
         10130 => x"2e",
         10131 => x"00",
         10132 => x"6f",
         10133 => x"65",
         10134 => x"75",
         10135 => x"64",
         10136 => x"61",
         10137 => x"74",
         10138 => x"6f",
         10139 => x"73",
         10140 => x"6d",
         10141 => x"64",
         10142 => x"00",
         10143 => x"74",
         10144 => x"20",
         10145 => x"6e",
         10146 => x"00",
         10147 => x"6e",
         10148 => x"2e",
         10149 => x"00",
         10150 => x"62",
         10151 => x"67",
         10152 => x"74",
         10153 => x"75",
         10154 => x"2e",
         10155 => x"00",
         10156 => x"25",
         10157 => x"64",
         10158 => x"3a",
         10159 => x"25",
         10160 => x"64",
         10161 => x"00",
         10162 => x"20",
         10163 => x"66",
         10164 => x"72",
         10165 => x"6f",
         10166 => x"00",
         10167 => x"72",
         10168 => x"53",
         10169 => x"63",
         10170 => x"69",
         10171 => x"00",
         10172 => x"65",
         10173 => x"65",
         10174 => x"6d",
         10175 => x"6d",
         10176 => x"65",
         10177 => x"00",
         10178 => x"20",
         10179 => x"53",
         10180 => x"4d",
         10181 => x"25",
         10182 => x"3a",
         10183 => x"58",
         10184 => x"00",
         10185 => x"20",
         10186 => x"41",
         10187 => x"20",
         10188 => x"25",
         10189 => x"3a",
         10190 => x"58",
         10191 => x"00",
         10192 => x"20",
         10193 => x"4e",
         10194 => x"41",
         10195 => x"25",
         10196 => x"3a",
         10197 => x"58",
         10198 => x"00",
         10199 => x"20",
         10200 => x"4d",
         10201 => x"20",
         10202 => x"25",
         10203 => x"3a",
         10204 => x"58",
         10205 => x"00",
         10206 => x"20",
         10207 => x"20",
         10208 => x"20",
         10209 => x"25",
         10210 => x"3a",
         10211 => x"58",
         10212 => x"00",
         10213 => x"20",
         10214 => x"43",
         10215 => x"20",
         10216 => x"44",
         10217 => x"63",
         10218 => x"3d",
         10219 => x"64",
         10220 => x"00",
         10221 => x"20",
         10222 => x"45",
         10223 => x"20",
         10224 => x"54",
         10225 => x"72",
         10226 => x"3d",
         10227 => x"64",
         10228 => x"00",
         10229 => x"20",
         10230 => x"52",
         10231 => x"52",
         10232 => x"43",
         10233 => x"6e",
         10234 => x"3d",
         10235 => x"64",
         10236 => x"00",
         10237 => x"20",
         10238 => x"48",
         10239 => x"45",
         10240 => x"53",
         10241 => x"00",
         10242 => x"20",
         10243 => x"49",
         10244 => x"00",
         10245 => x"20",
         10246 => x"54",
         10247 => x"00",
         10248 => x"20",
         10249 => x"00",
         10250 => x"20",
         10251 => x"00",
         10252 => x"72",
         10253 => x"65",
         10254 => x"00",
         10255 => x"20",
         10256 => x"20",
         10257 => x"65",
         10258 => x"65",
         10259 => x"72",
         10260 => x"64",
         10261 => x"73",
         10262 => x"25",
         10263 => x"0a",
         10264 => x"00",
         10265 => x"20",
         10266 => x"20",
         10267 => x"6f",
         10268 => x"53",
         10269 => x"74",
         10270 => x"64",
         10271 => x"73",
         10272 => x"25",
         10273 => x"0a",
         10274 => x"00",
         10275 => x"20",
         10276 => x"63",
         10277 => x"74",
         10278 => x"20",
         10279 => x"72",
         10280 => x"20",
         10281 => x"20",
         10282 => x"25",
         10283 => x"0a",
         10284 => x"00",
         10285 => x"63",
         10286 => x"00",
         10287 => x"20",
         10288 => x"20",
         10289 => x"20",
         10290 => x"20",
         10291 => x"20",
         10292 => x"20",
         10293 => x"20",
         10294 => x"25",
         10295 => x"0a",
         10296 => x"00",
         10297 => x"20",
         10298 => x"74",
         10299 => x"43",
         10300 => x"6b",
         10301 => x"65",
         10302 => x"20",
         10303 => x"20",
         10304 => x"25",
         10305 => x"30",
         10306 => x"48",
         10307 => x"00",
         10308 => x"20",
         10309 => x"41",
         10310 => x"6c",
         10311 => x"20",
         10312 => x"71",
         10313 => x"20",
         10314 => x"20",
         10315 => x"25",
         10316 => x"30",
         10317 => x"48",
         10318 => x"00",
         10319 => x"20",
         10320 => x"68",
         10321 => x"65",
         10322 => x"52",
         10323 => x"43",
         10324 => x"6b",
         10325 => x"65",
         10326 => x"25",
         10327 => x"30",
         10328 => x"48",
         10329 => x"00",
         10330 => x"6c",
         10331 => x"00",
         10332 => x"69",
         10333 => x"00",
         10334 => x"78",
         10335 => x"00",
         10336 => x"00",
         10337 => x"6d",
         10338 => x"00",
         10339 => x"6e",
         10340 => x"00",
         10341 => x"f0",
         10342 => x"00",
         10343 => x"02",
         10344 => x"ec",
         10345 => x"00",
         10346 => x"03",
         10347 => x"e8",
         10348 => x"00",
         10349 => x"04",
         10350 => x"e4",
         10351 => x"00",
         10352 => x"05",
         10353 => x"e0",
         10354 => x"00",
         10355 => x"06",
         10356 => x"dc",
         10357 => x"00",
         10358 => x"07",
         10359 => x"d8",
         10360 => x"00",
         10361 => x"01",
         10362 => x"d4",
         10363 => x"00",
         10364 => x"08",
         10365 => x"d0",
         10366 => x"00",
         10367 => x"0b",
         10368 => x"cc",
         10369 => x"00",
         10370 => x"09",
         10371 => x"c8",
         10372 => x"00",
         10373 => x"0a",
         10374 => x"c4",
         10375 => x"00",
         10376 => x"0d",
         10377 => x"c0",
         10378 => x"00",
         10379 => x"0c",
         10380 => x"bc",
         10381 => x"00",
         10382 => x"0e",
         10383 => x"b8",
         10384 => x"00",
         10385 => x"0f",
         10386 => x"b4",
         10387 => x"00",
         10388 => x"0f",
         10389 => x"b0",
         10390 => x"00",
         10391 => x"10",
         10392 => x"ac",
         10393 => x"00",
         10394 => x"11",
         10395 => x"a8",
         10396 => x"00",
         10397 => x"12",
         10398 => x"a4",
         10399 => x"00",
         10400 => x"13",
         10401 => x"a0",
         10402 => x"00",
         10403 => x"14",
         10404 => x"9c",
         10405 => x"00",
         10406 => x"15",
         10407 => x"00",
         10408 => x"00",
         10409 => x"00",
         10410 => x"00",
         10411 => x"7e",
         10412 => x"7e",
         10413 => x"7e",
         10414 => x"00",
         10415 => x"7e",
         10416 => x"7e",
         10417 => x"7e",
         10418 => x"00",
         10419 => x"00",
         10420 => x"00",
         10421 => x"00",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"74",
         10430 => x"00",
         10431 => x"74",
         10432 => x"00",
         10433 => x"00",
         10434 => x"6c",
         10435 => x"25",
         10436 => x"00",
         10437 => x"6c",
         10438 => x"74",
         10439 => x"65",
         10440 => x"20",
         10441 => x"20",
         10442 => x"74",
         10443 => x"20",
         10444 => x"65",
         10445 => x"20",
         10446 => x"2e",
         10447 => x"00",
         10448 => x"6e",
         10449 => x"6f",
         10450 => x"2f",
         10451 => x"61",
         10452 => x"68",
         10453 => x"6f",
         10454 => x"66",
         10455 => x"2c",
         10456 => x"73",
         10457 => x"69",
         10458 => x"00",
         10459 => x"00",
         10460 => x"3c",
         10461 => x"7f",
         10462 => x"00",
         10463 => x"3d",
         10464 => x"00",
         10465 => x"00",
         10466 => x"33",
         10467 => x"00",
         10468 => x"4d",
         10469 => x"53",
         10470 => x"00",
         10471 => x"4e",
         10472 => x"20",
         10473 => x"46",
         10474 => x"32",
         10475 => x"00",
         10476 => x"4e",
         10477 => x"20",
         10478 => x"46",
         10479 => x"20",
         10480 => x"00",
         10481 => x"6c",
         10482 => x"00",
         10483 => x"00",
         10484 => x"00",
         10485 => x"07",
         10486 => x"12",
         10487 => x"1c",
         10488 => x"00",
         10489 => x"41",
         10490 => x"80",
         10491 => x"49",
         10492 => x"8f",
         10493 => x"4f",
         10494 => x"55",
         10495 => x"9b",
         10496 => x"9f",
         10497 => x"55",
         10498 => x"a7",
         10499 => x"ab",
         10500 => x"af",
         10501 => x"b3",
         10502 => x"b7",
         10503 => x"bb",
         10504 => x"bf",
         10505 => x"c3",
         10506 => x"c7",
         10507 => x"cb",
         10508 => x"cf",
         10509 => x"d3",
         10510 => x"d7",
         10511 => x"db",
         10512 => x"df",
         10513 => x"e3",
         10514 => x"e7",
         10515 => x"eb",
         10516 => x"ef",
         10517 => x"f3",
         10518 => x"f7",
         10519 => x"fb",
         10520 => x"ff",
         10521 => x"3b",
         10522 => x"2f",
         10523 => x"3a",
         10524 => x"7c",
         10525 => x"00",
         10526 => x"04",
         10527 => x"40",
         10528 => x"00",
         10529 => x"00",
         10530 => x"02",
         10531 => x"08",
         10532 => x"20",
         10533 => x"00",
         10534 => x"fc",
         10535 => x"e2",
         10536 => x"e0",
         10537 => x"e7",
         10538 => x"eb",
         10539 => x"ef",
         10540 => x"ec",
         10541 => x"c5",
         10542 => x"e6",
         10543 => x"f4",
         10544 => x"f2",
         10545 => x"f9",
         10546 => x"d6",
         10547 => x"a2",
         10548 => x"a5",
         10549 => x"92",
         10550 => x"ed",
         10551 => x"fa",
         10552 => x"d1",
         10553 => x"ba",
         10554 => x"10",
         10555 => x"bd",
         10556 => x"a1",
         10557 => x"bb",
         10558 => x"92",
         10559 => x"02",
         10560 => x"61",
         10561 => x"56",
         10562 => x"63",
         10563 => x"57",
         10564 => x"5c",
         10565 => x"10",
         10566 => x"34",
         10567 => x"1c",
         10568 => x"3c",
         10569 => x"5f",
         10570 => x"54",
         10571 => x"66",
         10572 => x"50",
         10573 => x"67",
         10574 => x"64",
         10575 => x"59",
         10576 => x"52",
         10577 => x"6b",
         10578 => x"18",
         10579 => x"88",
         10580 => x"8c",
         10581 => x"80",
         10582 => x"df",
         10583 => x"c0",
         10584 => x"c3",
         10585 => x"c4",
         10586 => x"98",
         10587 => x"b4",
         10588 => x"c6",
         10589 => x"29",
         10590 => x"b1",
         10591 => x"64",
         10592 => x"21",
         10593 => x"48",
         10594 => x"19",
         10595 => x"1a",
         10596 => x"b2",
         10597 => x"a0",
         10598 => x"1a",
         10599 => x"17",
         10600 => x"07",
         10601 => x"01",
         10602 => x"00",
         10603 => x"32",
         10604 => x"39",
         10605 => x"4a",
         10606 => x"79",
         10607 => x"80",
         10608 => x"43",
         10609 => x"82",
         10610 => x"84",
         10611 => x"86",
         10612 => x"87",
         10613 => x"8a",
         10614 => x"8b",
         10615 => x"8e",
         10616 => x"90",
         10617 => x"91",
         10618 => x"94",
         10619 => x"96",
         10620 => x"98",
         10621 => x"3d",
         10622 => x"9c",
         10623 => x"20",
         10624 => x"a0",
         10625 => x"a2",
         10626 => x"a4",
         10627 => x"a6",
         10628 => x"a7",
         10629 => x"aa",
         10630 => x"ac",
         10631 => x"ae",
         10632 => x"af",
         10633 => x"b2",
         10634 => x"b3",
         10635 => x"b5",
         10636 => x"b8",
         10637 => x"ba",
         10638 => x"bc",
         10639 => x"be",
         10640 => x"c0",
         10641 => x"c2",
         10642 => x"c4",
         10643 => x"c4",
         10644 => x"c8",
         10645 => x"ca",
         10646 => x"ca",
         10647 => x"10",
         10648 => x"01",
         10649 => x"de",
         10650 => x"f3",
         10651 => x"f1",
         10652 => x"f4",
         10653 => x"28",
         10654 => x"12",
         10655 => x"09",
         10656 => x"3b",
         10657 => x"3d",
         10658 => x"3f",
         10659 => x"41",
         10660 => x"46",
         10661 => x"53",
         10662 => x"81",
         10663 => x"55",
         10664 => x"8a",
         10665 => x"8f",
         10666 => x"90",
         10667 => x"5d",
         10668 => x"5f",
         10669 => x"61",
         10670 => x"94",
         10671 => x"65",
         10672 => x"67",
         10673 => x"96",
         10674 => x"62",
         10675 => x"6d",
         10676 => x"9c",
         10677 => x"71",
         10678 => x"73",
         10679 => x"9f",
         10680 => x"77",
         10681 => x"79",
         10682 => x"7b",
         10683 => x"64",
         10684 => x"7f",
         10685 => x"81",
         10686 => x"a9",
         10687 => x"85",
         10688 => x"87",
         10689 => x"44",
         10690 => x"b2",
         10691 => x"8d",
         10692 => x"8f",
         10693 => x"91",
         10694 => x"7b",
         10695 => x"fd",
         10696 => x"ff",
         10697 => x"04",
         10698 => x"88",
         10699 => x"8a",
         10700 => x"11",
         10701 => x"02",
         10702 => x"a3",
         10703 => x"08",
         10704 => x"03",
         10705 => x"8e",
         10706 => x"d8",
         10707 => x"f2",
         10708 => x"f9",
         10709 => x"f4",
         10710 => x"f6",
         10711 => x"f7",
         10712 => x"fa",
         10713 => x"30",
         10714 => x"50",
         10715 => x"60",
         10716 => x"8a",
         10717 => x"c1",
         10718 => x"cf",
         10719 => x"c0",
         10720 => x"44",
         10721 => x"26",
         10722 => x"00",
         10723 => x"01",
         10724 => x"00",
         10725 => x"a0",
         10726 => x"00",
         10727 => x"10",
         10728 => x"20",
         10729 => x"30",
         10730 => x"40",
         10731 => x"51",
         10732 => x"59",
         10733 => x"5b",
         10734 => x"5d",
         10735 => x"5f",
         10736 => x"08",
         10737 => x"0e",
         10738 => x"bb",
         10739 => x"c9",
         10740 => x"cb",
         10741 => x"db",
         10742 => x"f9",
         10743 => x"eb",
         10744 => x"fb",
         10745 => x"08",
         10746 => x"08",
         10747 => x"08",
         10748 => x"04",
         10749 => x"b9",
         10750 => x"bc",
         10751 => x"01",
         10752 => x"d0",
         10753 => x"e0",
         10754 => x"e5",
         10755 => x"ec",
         10756 => x"01",
         10757 => x"4e",
         10758 => x"32",
         10759 => x"10",
         10760 => x"01",
         10761 => x"d0",
         10762 => x"30",
         10763 => x"60",
         10764 => x"67",
         10765 => x"75",
         10766 => x"80",
         10767 => x"00",
         10768 => x"41",
         10769 => x"00",
         10770 => x"00",
         10771 => x"a0",
         10772 => x"00",
         10773 => x"00",
         10774 => x"00",
         10775 => x"a8",
         10776 => x"00",
         10777 => x"00",
         10778 => x"00",
         10779 => x"b0",
         10780 => x"00",
         10781 => x"00",
         10782 => x"00",
         10783 => x"b8",
         10784 => x"00",
         10785 => x"00",
         10786 => x"00",
         10787 => x"c0",
         10788 => x"00",
         10789 => x"00",
         10790 => x"00",
         10791 => x"c8",
         10792 => x"00",
         10793 => x"00",
         10794 => x"00",
         10795 => x"d0",
         10796 => x"00",
         10797 => x"00",
         10798 => x"00",
         10799 => x"d8",
         10800 => x"00",
         10801 => x"00",
         10802 => x"00",
         10803 => x"e0",
         10804 => x"00",
         10805 => x"00",
         10806 => x"00",
         10807 => x"e8",
         10808 => x"00",
         10809 => x"00",
         10810 => x"00",
         10811 => x"ec",
         10812 => x"00",
         10813 => x"00",
         10814 => x"00",
         10815 => x"f0",
         10816 => x"00",
         10817 => x"00",
         10818 => x"00",
         10819 => x"f4",
         10820 => x"00",
         10821 => x"00",
         10822 => x"00",
         10823 => x"f8",
         10824 => x"00",
         10825 => x"00",
         10826 => x"00",
         10827 => x"fc",
         10828 => x"00",
         10829 => x"00",
         10830 => x"00",
         10831 => x"00",
         10832 => x"00",
         10833 => x"00",
         10834 => x"00",
         10835 => x"04",
         10836 => x"00",
         10837 => x"00",
         10838 => x"00",
         10839 => x"0c",
         10840 => x"00",
         10841 => x"00",
         10842 => x"00",
         10843 => x"10",
         10844 => x"00",
         10845 => x"00",
         10846 => x"00",
         10847 => x"18",
         10848 => x"00",
         10849 => x"00",
         10850 => x"00",
         10851 => x"20",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"28",
         10856 => x"00",
         10857 => x"00",
         10858 => x"00",
         10859 => x"30",
         10860 => x"00",
         10861 => x"00",
         10862 => x"00",
         10863 => x"38",
         10864 => x"00",
         10865 => x"00",
         10866 => x"00",
         10867 => x"40",
         10868 => x"00",
         10869 => x"00",
         10870 => x"00",
         10871 => x"48",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"ff",
         10878 => x"00",
         10879 => x"ff",
         10880 => x"00",
         10881 => x"ff",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"ff",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"01",
         10895 => x"01",
         10896 => x"01",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"f4",
         10923 => x"00",
         10924 => x"fc",
         10925 => x"00",
         10926 => x"04",
         10927 => x"00",
         10928 => x"f3",
         10929 => x"f7",
         10930 => x"fb",
         10931 => x"ff",
         10932 => x"c3",
         10933 => x"e2",
         10934 => x"e6",
         10935 => x"f4",
         10936 => x"63",
         10937 => x"67",
         10938 => x"6a",
         10939 => x"2d",
         10940 => x"23",
         10941 => x"27",
         10942 => x"2c",
         10943 => x"49",
         10944 => x"03",
         10945 => x"07",
         10946 => x"0b",
         10947 => x"0f",
         10948 => x"13",
         10949 => x"17",
         10950 => x"52",
         10951 => x"3c",
         10952 => x"83",
         10953 => x"87",
         10954 => x"8b",
         10955 => x"8f",
         10956 => x"93",
         10957 => x"97",
         10958 => x"bc",
         10959 => x"c0",
         10960 => x"00",
         10961 => x"00",
         10962 => x"00",
         10963 => x"00",
         10964 => x"00",
         10965 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"d6",
           386 => x"f7",
           387 => x"d6",
           388 => x"80",
           389 => x"d6",
           390 => x"b2",
           391 => x"e4",
           392 => x"90",
           393 => x"e4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"84",
           400 => x"82",
           401 => x"94",
           402 => x"d6",
           403 => x"80",
           404 => x"d6",
           405 => x"c2",
           406 => x"e4",
           407 => x"90",
           408 => x"e4",
           409 => x"f7",
           410 => x"e4",
           411 => x"90",
           412 => x"e4",
           413 => x"a6",
           414 => x"e4",
           415 => x"90",
           416 => x"e4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"84",
           423 => x"82",
           424 => x"97",
           425 => x"d6",
           426 => x"80",
           427 => x"d6",
           428 => x"f9",
           429 => x"d6",
           430 => x"80",
           431 => x"d6",
           432 => x"fa",
           433 => x"d6",
           434 => x"80",
           435 => x"d6",
           436 => x"f3",
           437 => x"d6",
           438 => x"80",
           439 => x"d6",
           440 => x"f5",
           441 => x"d6",
           442 => x"80",
           443 => x"d6",
           444 => x"f6",
           445 => x"d6",
           446 => x"80",
           447 => x"d6",
           448 => x"ec",
           449 => x"d6",
           450 => x"80",
           451 => x"d6",
           452 => x"f9",
           453 => x"d6",
           454 => x"80",
           455 => x"d6",
           456 => x"f1",
           457 => x"d6",
           458 => x"80",
           459 => x"d6",
           460 => x"f4",
           461 => x"d6",
           462 => x"80",
           463 => x"d6",
           464 => x"fe",
           465 => x"d6",
           466 => x"80",
           467 => x"d6",
           468 => x"87",
           469 => x"d6",
           470 => x"80",
           471 => x"d6",
           472 => x"f8",
           473 => x"d6",
           474 => x"80",
           475 => x"d6",
           476 => x"82",
           477 => x"d6",
           478 => x"80",
           479 => x"d6",
           480 => x"83",
           481 => x"d6",
           482 => x"80",
           483 => x"d6",
           484 => x"83",
           485 => x"d6",
           486 => x"80",
           487 => x"d6",
           488 => x"8b",
           489 => x"d6",
           490 => x"80",
           491 => x"d6",
           492 => x"89",
           493 => x"d6",
           494 => x"80",
           495 => x"d6",
           496 => x"8e",
           497 => x"d6",
           498 => x"80",
           499 => x"d6",
           500 => x"84",
           501 => x"d6",
           502 => x"80",
           503 => x"d6",
           504 => x"91",
           505 => x"d6",
           506 => x"80",
           507 => x"d6",
           508 => x"92",
           509 => x"d6",
           510 => x"80",
           511 => x"d6",
           512 => x"fa",
           513 => x"d6",
           514 => x"80",
           515 => x"d6",
           516 => x"f9",
           517 => x"d6",
           518 => x"80",
           519 => x"d6",
           520 => x"fb",
           521 => x"d6",
           522 => x"80",
           523 => x"d6",
           524 => x"85",
           525 => x"d6",
           526 => x"80",
           527 => x"d6",
           528 => x"93",
           529 => x"d6",
           530 => x"80",
           531 => x"d6",
           532 => x"95",
           533 => x"d6",
           534 => x"80",
           535 => x"d6",
           536 => x"98",
           537 => x"d6",
           538 => x"80",
           539 => x"d6",
           540 => x"eb",
           541 => x"d6",
           542 => x"80",
           543 => x"d6",
           544 => x"9b",
           545 => x"d6",
           546 => x"80",
           547 => x"d6",
           548 => x"a9",
           549 => x"d6",
           550 => x"80",
           551 => x"d6",
           552 => x"a7",
           553 => x"d6",
           554 => x"80",
           555 => x"d6",
           556 => x"ab",
           557 => x"d6",
           558 => x"80",
           559 => x"d6",
           560 => x"ad",
           561 => x"d6",
           562 => x"80",
           563 => x"d6",
           564 => x"af",
           565 => x"d6",
           566 => x"80",
           567 => x"d6",
           568 => x"f3",
           569 => x"d6",
           570 => x"80",
           571 => x"d6",
           572 => x"f4",
           573 => x"d6",
           574 => x"80",
           575 => x"d6",
           576 => x"f8",
           577 => x"d6",
           578 => x"80",
           579 => x"d6",
           580 => x"d7",
           581 => x"d6",
           582 => x"80",
           583 => x"d6",
           584 => x"a5",
           585 => x"d6",
           586 => x"80",
           587 => x"d6",
           588 => x"a6",
           589 => x"d6",
           590 => x"80",
           591 => x"d6",
           592 => x"aa",
           593 => x"d6",
           594 => x"80",
           595 => x"d6",
           596 => x"a2",
           597 => x"d6",
           598 => x"80",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"d6",
           623 => x"f2",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"e4",
           631 => x"d6",
           632 => x"3d",
           633 => x"e4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"e4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"e4",
           651 => x"d6",
           652 => x"82",
           653 => x"fb",
           654 => x"d6",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"e4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"e4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"d6",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"d6",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"e4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"e4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"e4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"d6",
           712 => x"05",
           713 => x"d6",
           714 => x"05",
           715 => x"d6",
           716 => x"05",
           717 => x"d8",
           718 => x"0d",
           719 => x"0c",
           720 => x"e4",
           721 => x"d6",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"d6",
           726 => x"05",
           727 => x"e4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"d6",
           732 => x"05",
           733 => x"e4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"d8",
           743 => x"d6",
           744 => x"05",
           745 => x"e4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"e4",
           751 => x"08",
           752 => x"d8",
           753 => x"3d",
           754 => x"e4",
           755 => x"d6",
           756 => x"82",
           757 => x"fb",
           758 => x"d6",
           759 => x"05",
           760 => x"e4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"e4",
           778 => x"d6",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"d6",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"d6",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"d6",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"d6",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"d6",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"e4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"e4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"e4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"d6",
           848 => x"05",
           849 => x"e4",
           850 => x"33",
           851 => x"e4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"d6",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"d6",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"e4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"d6",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"d6",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"ae",
           901 => x"08",
           902 => x"53",
           903 => x"d6",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"d6",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"e4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"e4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"e4",
           927 => x"22",
           928 => x"51",
           929 => x"d6",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"e4",
           935 => x"22",
           936 => x"51",
           937 => x"d6",
           938 => x"05",
           939 => x"39",
           940 => x"d6",
           941 => x"05",
           942 => x"e4",
           943 => x"22",
           944 => x"53",
           945 => x"e4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"e4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"e4",
           955 => x"0c",
           956 => x"53",
           957 => x"e4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"d6",
           965 => x"05",
           966 => x"e4",
           967 => x"08",
           968 => x"d6",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"d6",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"e4",
           987 => x"23",
           988 => x"d6",
           989 => x"05",
           990 => x"8a",
           991 => x"d8",
           992 => x"82",
           993 => x"f4",
           994 => x"d6",
           995 => x"05",
           996 => x"d6",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"e4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"e4",
          1007 => x"0c",
          1008 => x"d6",
          1009 => x"05",
          1010 => x"e4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"d6",
          1020 => x"05",
          1021 => x"a2",
          1022 => x"d6",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"e4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"d6",
          1031 => x"05",
          1032 => x"e4",
          1033 => x"22",
          1034 => x"e4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"d6",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"e4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"e4",
          1050 => x"0c",
          1051 => x"d6",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"e4",
          1061 => x"0c",
          1062 => x"e4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"d6",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"d6",
          1074 => x"05",
          1075 => x"d6",
          1076 => x"05",
          1077 => x"e4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"d6",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"e4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"e4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"e4",
          1106 => x"0c",
          1107 => x"d6",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"e4",
          1117 => x"0c",
          1118 => x"e4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"d6",
          1130 => x"05",
          1131 => x"e4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"9e",
          1137 => x"d8",
          1138 => x"75",
          1139 => x"e4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"d6",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"e4",
          1154 => x"34",
          1155 => x"d6",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"e4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"e4",
          1166 => x"08",
          1167 => x"d6",
          1168 => x"05",
          1169 => x"e4",
          1170 => x"22",
          1171 => x"d6",
          1172 => x"05",
          1173 => x"a3",
          1174 => x"d6",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"e4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"d6",
          1187 => x"05",
          1188 => x"e4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"d6",
          1193 => x"05",
          1194 => x"51",
          1195 => x"d6",
          1196 => x"05",
          1197 => x"e4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"e4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"e4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"e4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"e4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"d6",
          1227 => x"05",
          1228 => x"e4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"e4",
          1245 => x"23",
          1246 => x"d6",
          1247 => x"05",
          1248 => x"d6",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"d6",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"e4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"d6",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"e4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"d6",
          1281 => x"05",
          1282 => x"e4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"e4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"e4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"e4",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"e4",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"e4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"d6",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"e4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"d6",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"e4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"e4",
          1338 => x"08",
          1339 => x"e4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"e4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"e4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"e4",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"e4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"e4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"e4",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"d6",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"e4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"d6",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"e4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"d6",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"e4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"d6",
          1452 => x"05",
          1453 => x"d6",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"d6",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"d6",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"d6",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"e4",
          1494 => x"23",
          1495 => x"d6",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"e4",
          1501 => x"08",
          1502 => x"e4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"d6",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"d6",
          1513 => x"3d",
          1514 => x"e4",
          1515 => x"d6",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"f2",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"d6",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"e4",
          1531 => x"0d",
          1532 => x"d6",
          1533 => x"05",
          1534 => x"bc",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"e4",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"e4",
          1547 => x"08",
          1548 => x"d6",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"e4",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"e4",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"d8",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"e4",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"d6",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"e4",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"e4",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"e4",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"d6",
          1612 => x"05",
          1613 => x"e4",
          1614 => x"08",
          1615 => x"e4",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"e4",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"d6",
          1631 => x"3d",
          1632 => x"e4",
          1633 => x"d6",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"f2",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"d8",
          1641 => x"d6",
          1642 => x"84",
          1643 => x"d6",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"d6",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"d6",
          1665 => x"05",
          1666 => x"e4",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"e4",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"e4",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"d6",
          1702 => x"05",
          1703 => x"d6",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"d6",
          1709 => x"05",
          1710 => x"d8",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"e4",
          1714 => x"d6",
          1715 => x"3d",
          1716 => x"e4",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"d6",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"e4",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"d6",
          1756 => x"05",
          1757 => x"70",
          1758 => x"e4",
          1759 => x"0c",
          1760 => x"d6",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"d6",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"e4",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"d6",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"d6",
          1791 => x"05",
          1792 => x"e4",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"e4",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"e4",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"e4",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"e4",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"d6",
          1838 => x"05",
          1839 => x"e4",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"d6",
          1849 => x"05",
          1850 => x"e4",
          1851 => x"08",
          1852 => x"d6",
          1853 => x"05",
          1854 => x"81",
          1855 => x"d6",
          1856 => x"05",
          1857 => x"e4",
          1858 => x"08",
          1859 => x"e4",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"d6",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"d6",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"d6",
          1875 => x"05",
          1876 => x"81",
          1877 => x"d6",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"d6",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"d6",
          1886 => x"05",
          1887 => x"e4",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"e4",
          1892 => x"08",
          1893 => x"d6",
          1894 => x"05",
          1895 => x"e4",
          1896 => x"08",
          1897 => x"d6",
          1898 => x"05",
          1899 => x"e4",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"d6",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"d6",
          1909 => x"05",
          1910 => x"71",
          1911 => x"d6",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"e4",
          1917 => x"08",
          1918 => x"d8",
          1919 => x"3d",
          1920 => x"e4",
          1921 => x"d6",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"d6",
          1925 => x"05",
          1926 => x"e4",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"d6",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"d6",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"e4",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"d6",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"e4",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"e4",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"e4",
          1973 => x"08",
          1974 => x"d8",
          1975 => x"3d",
          1976 => x"e4",
          1977 => x"d6",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"d6",
          1981 => x"05",
          1982 => x"e4",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"d6",
          1988 => x"05",
          1989 => x"80",
          1990 => x"d6",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"d6",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"d6",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"e4",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"d6",
          2016 => x"05",
          2017 => x"d6",
          2018 => x"85",
          2019 => x"d6",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"e4",
          2030 => x"08",
          2031 => x"d6",
          2032 => x"05",
          2033 => x"e4",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"d6",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"e4",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"e4",
          2052 => x"08",
          2053 => x"d6",
          2054 => x"05",
          2055 => x"e4",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"e4",
          2069 => x"08",
          2070 => x"d6",
          2071 => x"05",
          2072 => x"e4",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"e4",
          2077 => x"0c",
          2078 => x"d6",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"d6",
          2092 => x"3d",
          2093 => x"e4",
          2094 => x"d6",
          2095 => x"82",
          2096 => x"fa",
          2097 => x"d6",
          2098 => x"05",
          2099 => x"d6",
          2100 => x"05",
          2101 => x"8d",
          2102 => x"d8",
          2103 => x"d6",
          2104 => x"05",
          2105 => x"e4",
          2106 => x"08",
          2107 => x"53",
          2108 => x"e3",
          2109 => x"d6",
          2110 => x"82",
          2111 => x"fc",
          2112 => x"82",
          2113 => x"fc",
          2114 => x"38",
          2115 => x"d6",
          2116 => x"05",
          2117 => x"82",
          2118 => x"fc",
          2119 => x"d6",
          2120 => x"05",
          2121 => x"80",
          2122 => x"d6",
          2123 => x"05",
          2124 => x"d6",
          2125 => x"05",
          2126 => x"d6",
          2127 => x"05",
          2128 => x"a2",
          2129 => x"d8",
          2130 => x"d6",
          2131 => x"05",
          2132 => x"d6",
          2133 => x"05",
          2134 => x"d8",
          2135 => x"0d",
          2136 => x"0c",
          2137 => x"e4",
          2138 => x"d6",
          2139 => x"3d",
          2140 => x"e4",
          2141 => x"08",
          2142 => x"08",
          2143 => x"82",
          2144 => x"8c",
          2145 => x"38",
          2146 => x"d6",
          2147 => x"05",
          2148 => x"39",
          2149 => x"08",
          2150 => x"52",
          2151 => x"d6",
          2152 => x"05",
          2153 => x"82",
          2154 => x"f8",
          2155 => x"81",
          2156 => x"51",
          2157 => x"9f",
          2158 => x"e4",
          2159 => x"08",
          2160 => x"d6",
          2161 => x"05",
          2162 => x"e4",
          2163 => x"08",
          2164 => x"38",
          2165 => x"82",
          2166 => x"f8",
          2167 => x"05",
          2168 => x"08",
          2169 => x"82",
          2170 => x"f8",
          2171 => x"d6",
          2172 => x"05",
          2173 => x"82",
          2174 => x"fc",
          2175 => x"82",
          2176 => x"fc",
          2177 => x"d6",
          2178 => x"3d",
          2179 => x"e4",
          2180 => x"d6",
          2181 => x"82",
          2182 => x"fe",
          2183 => x"d6",
          2184 => x"05",
          2185 => x"e4",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"80",
          2189 => x"38",
          2190 => x"08",
          2191 => x"81",
          2192 => x"e4",
          2193 => x"0c",
          2194 => x"08",
          2195 => x"ff",
          2196 => x"e4",
          2197 => x"0c",
          2198 => x"08",
          2199 => x"80",
          2200 => x"82",
          2201 => x"8c",
          2202 => x"70",
          2203 => x"08",
          2204 => x"52",
          2205 => x"34",
          2206 => x"08",
          2207 => x"81",
          2208 => x"e4",
          2209 => x"0c",
          2210 => x"82",
          2211 => x"88",
          2212 => x"82",
          2213 => x"51",
          2214 => x"82",
          2215 => x"04",
          2216 => x"08",
          2217 => x"e4",
          2218 => x"0d",
          2219 => x"d6",
          2220 => x"05",
          2221 => x"e4",
          2222 => x"08",
          2223 => x"38",
          2224 => x"08",
          2225 => x"30",
          2226 => x"08",
          2227 => x"80",
          2228 => x"e4",
          2229 => x"0c",
          2230 => x"08",
          2231 => x"8a",
          2232 => x"82",
          2233 => x"f4",
          2234 => x"d6",
          2235 => x"05",
          2236 => x"e4",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"8c",
          2242 => x"82",
          2243 => x"8c",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"fc",
          2248 => x"38",
          2249 => x"d6",
          2250 => x"05",
          2251 => x"e4",
          2252 => x"08",
          2253 => x"08",
          2254 => x"80",
          2255 => x"e4",
          2256 => x"08",
          2257 => x"e4",
          2258 => x"08",
          2259 => x"3f",
          2260 => x"08",
          2261 => x"e4",
          2262 => x"0c",
          2263 => x"e4",
          2264 => x"08",
          2265 => x"38",
          2266 => x"08",
          2267 => x"30",
          2268 => x"08",
          2269 => x"82",
          2270 => x"f8",
          2271 => x"82",
          2272 => x"54",
          2273 => x"82",
          2274 => x"04",
          2275 => x"08",
          2276 => x"e4",
          2277 => x"0d",
          2278 => x"d6",
          2279 => x"05",
          2280 => x"e4",
          2281 => x"08",
          2282 => x"38",
          2283 => x"08",
          2284 => x"30",
          2285 => x"08",
          2286 => x"81",
          2287 => x"e4",
          2288 => x"0c",
          2289 => x"08",
          2290 => x"80",
          2291 => x"82",
          2292 => x"8c",
          2293 => x"82",
          2294 => x"8c",
          2295 => x"53",
          2296 => x"08",
          2297 => x"52",
          2298 => x"08",
          2299 => x"51",
          2300 => x"82",
          2301 => x"70",
          2302 => x"08",
          2303 => x"54",
          2304 => x"08",
          2305 => x"80",
          2306 => x"82",
          2307 => x"f8",
          2308 => x"82",
          2309 => x"f8",
          2310 => x"d6",
          2311 => x"05",
          2312 => x"d6",
          2313 => x"87",
          2314 => x"d6",
          2315 => x"82",
          2316 => x"02",
          2317 => x"0c",
          2318 => x"80",
          2319 => x"e4",
          2320 => x"08",
          2321 => x"e4",
          2322 => x"08",
          2323 => x"3f",
          2324 => x"08",
          2325 => x"d8",
          2326 => x"3d",
          2327 => x"e4",
          2328 => x"d6",
          2329 => x"82",
          2330 => x"fd",
          2331 => x"53",
          2332 => x"08",
          2333 => x"52",
          2334 => x"08",
          2335 => x"51",
          2336 => x"d6",
          2337 => x"82",
          2338 => x"54",
          2339 => x"82",
          2340 => x"04",
          2341 => x"08",
          2342 => x"e4",
          2343 => x"0d",
          2344 => x"d6",
          2345 => x"05",
          2346 => x"82",
          2347 => x"f8",
          2348 => x"d6",
          2349 => x"05",
          2350 => x"e4",
          2351 => x"08",
          2352 => x"82",
          2353 => x"fc",
          2354 => x"2e",
          2355 => x"0b",
          2356 => x"08",
          2357 => x"24",
          2358 => x"d6",
          2359 => x"05",
          2360 => x"d6",
          2361 => x"05",
          2362 => x"e4",
          2363 => x"08",
          2364 => x"e4",
          2365 => x"0c",
          2366 => x"82",
          2367 => x"fc",
          2368 => x"2e",
          2369 => x"82",
          2370 => x"8c",
          2371 => x"d6",
          2372 => x"05",
          2373 => x"38",
          2374 => x"08",
          2375 => x"82",
          2376 => x"8c",
          2377 => x"82",
          2378 => x"88",
          2379 => x"d6",
          2380 => x"05",
          2381 => x"e4",
          2382 => x"08",
          2383 => x"e4",
          2384 => x"0c",
          2385 => x"08",
          2386 => x"81",
          2387 => x"e4",
          2388 => x"0c",
          2389 => x"08",
          2390 => x"81",
          2391 => x"e4",
          2392 => x"0c",
          2393 => x"82",
          2394 => x"90",
          2395 => x"2e",
          2396 => x"d6",
          2397 => x"05",
          2398 => x"d6",
          2399 => x"05",
          2400 => x"39",
          2401 => x"08",
          2402 => x"70",
          2403 => x"08",
          2404 => x"51",
          2405 => x"08",
          2406 => x"82",
          2407 => x"85",
          2408 => x"d6",
          2409 => x"82",
          2410 => x"02",
          2411 => x"0c",
          2412 => x"80",
          2413 => x"e4",
          2414 => x"34",
          2415 => x"08",
          2416 => x"53",
          2417 => x"82",
          2418 => x"88",
          2419 => x"08",
          2420 => x"33",
          2421 => x"d6",
          2422 => x"05",
          2423 => x"ff",
          2424 => x"a0",
          2425 => x"06",
          2426 => x"d6",
          2427 => x"05",
          2428 => x"81",
          2429 => x"53",
          2430 => x"d6",
          2431 => x"05",
          2432 => x"ad",
          2433 => x"06",
          2434 => x"0b",
          2435 => x"08",
          2436 => x"82",
          2437 => x"88",
          2438 => x"08",
          2439 => x"0c",
          2440 => x"53",
          2441 => x"d6",
          2442 => x"05",
          2443 => x"e4",
          2444 => x"33",
          2445 => x"2e",
          2446 => x"81",
          2447 => x"d6",
          2448 => x"05",
          2449 => x"81",
          2450 => x"70",
          2451 => x"72",
          2452 => x"e4",
          2453 => x"34",
          2454 => x"08",
          2455 => x"82",
          2456 => x"e8",
          2457 => x"d6",
          2458 => x"05",
          2459 => x"2e",
          2460 => x"d6",
          2461 => x"05",
          2462 => x"2e",
          2463 => x"cd",
          2464 => x"82",
          2465 => x"f4",
          2466 => x"d6",
          2467 => x"05",
          2468 => x"81",
          2469 => x"70",
          2470 => x"72",
          2471 => x"e4",
          2472 => x"34",
          2473 => x"82",
          2474 => x"e4",
          2475 => x"34",
          2476 => x"08",
          2477 => x"70",
          2478 => x"71",
          2479 => x"51",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"fe",
          2483 => x"e4",
          2484 => x"33",
          2485 => x"26",
          2486 => x"0b",
          2487 => x"08",
          2488 => x"83",
          2489 => x"d6",
          2490 => x"05",
          2491 => x"73",
          2492 => x"82",
          2493 => x"f8",
          2494 => x"72",
          2495 => x"38",
          2496 => x"0b",
          2497 => x"08",
          2498 => x"82",
          2499 => x"0b",
          2500 => x"08",
          2501 => x"b2",
          2502 => x"e4",
          2503 => x"33",
          2504 => x"27",
          2505 => x"d6",
          2506 => x"05",
          2507 => x"b9",
          2508 => x"8d",
          2509 => x"82",
          2510 => x"ec",
          2511 => x"a5",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"0b",
          2515 => x"08",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"a0",
          2519 => x"cf",
          2520 => x"e4",
          2521 => x"33",
          2522 => x"73",
          2523 => x"82",
          2524 => x"f8",
          2525 => x"11",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"d6",
          2529 => x"05",
          2530 => x"51",
          2531 => x"d6",
          2532 => x"05",
          2533 => x"e4",
          2534 => x"33",
          2535 => x"27",
          2536 => x"d6",
          2537 => x"05",
          2538 => x"51",
          2539 => x"d6",
          2540 => x"05",
          2541 => x"e4",
          2542 => x"33",
          2543 => x"26",
          2544 => x"0b",
          2545 => x"08",
          2546 => x"81",
          2547 => x"d6",
          2548 => x"05",
          2549 => x"e4",
          2550 => x"33",
          2551 => x"74",
          2552 => x"80",
          2553 => x"e4",
          2554 => x"0c",
          2555 => x"82",
          2556 => x"f4",
          2557 => x"82",
          2558 => x"fc",
          2559 => x"82",
          2560 => x"f8",
          2561 => x"12",
          2562 => x"08",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"51",
          2568 => x"72",
          2569 => x"e4",
          2570 => x"34",
          2571 => x"82",
          2572 => x"f0",
          2573 => x"72",
          2574 => x"38",
          2575 => x"08",
          2576 => x"30",
          2577 => x"08",
          2578 => x"82",
          2579 => x"8c",
          2580 => x"d6",
          2581 => x"05",
          2582 => x"53",
          2583 => x"d6",
          2584 => x"05",
          2585 => x"e4",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"82",
          2589 => x"04",
          2590 => x"08",
          2591 => x"e4",
          2592 => x"0d",
          2593 => x"d6",
          2594 => x"05",
          2595 => x"e4",
          2596 => x"08",
          2597 => x"0c",
          2598 => x"08",
          2599 => x"70",
          2600 => x"72",
          2601 => x"82",
          2602 => x"f8",
          2603 => x"81",
          2604 => x"72",
          2605 => x"81",
          2606 => x"82",
          2607 => x"88",
          2608 => x"08",
          2609 => x"0c",
          2610 => x"82",
          2611 => x"f8",
          2612 => x"72",
          2613 => x"81",
          2614 => x"81",
          2615 => x"e4",
          2616 => x"34",
          2617 => x"08",
          2618 => x"70",
          2619 => x"71",
          2620 => x"51",
          2621 => x"82",
          2622 => x"f8",
          2623 => x"d6",
          2624 => x"05",
          2625 => x"b0",
          2626 => x"06",
          2627 => x"82",
          2628 => x"88",
          2629 => x"08",
          2630 => x"0c",
          2631 => x"53",
          2632 => x"d6",
          2633 => x"05",
          2634 => x"e4",
          2635 => x"33",
          2636 => x"08",
          2637 => x"82",
          2638 => x"e8",
          2639 => x"e2",
          2640 => x"82",
          2641 => x"e8",
          2642 => x"f8",
          2643 => x"80",
          2644 => x"0b",
          2645 => x"08",
          2646 => x"82",
          2647 => x"88",
          2648 => x"08",
          2649 => x"0c",
          2650 => x"53",
          2651 => x"d6",
          2652 => x"05",
          2653 => x"39",
          2654 => x"d6",
          2655 => x"05",
          2656 => x"e4",
          2657 => x"08",
          2658 => x"05",
          2659 => x"08",
          2660 => x"33",
          2661 => x"08",
          2662 => x"80",
          2663 => x"d6",
          2664 => x"05",
          2665 => x"a0",
          2666 => x"81",
          2667 => x"e4",
          2668 => x"0c",
          2669 => x"82",
          2670 => x"f8",
          2671 => x"af",
          2672 => x"38",
          2673 => x"08",
          2674 => x"53",
          2675 => x"83",
          2676 => x"80",
          2677 => x"e4",
          2678 => x"0c",
          2679 => x"88",
          2680 => x"e4",
          2681 => x"34",
          2682 => x"d6",
          2683 => x"05",
          2684 => x"73",
          2685 => x"82",
          2686 => x"f8",
          2687 => x"72",
          2688 => x"38",
          2689 => x"0b",
          2690 => x"08",
          2691 => x"82",
          2692 => x"0b",
          2693 => x"08",
          2694 => x"80",
          2695 => x"e4",
          2696 => x"0c",
          2697 => x"08",
          2698 => x"53",
          2699 => x"81",
          2700 => x"d6",
          2701 => x"05",
          2702 => x"e0",
          2703 => x"38",
          2704 => x"08",
          2705 => x"e0",
          2706 => x"72",
          2707 => x"08",
          2708 => x"82",
          2709 => x"f8",
          2710 => x"11",
          2711 => x"82",
          2712 => x"f8",
          2713 => x"d6",
          2714 => x"05",
          2715 => x"73",
          2716 => x"82",
          2717 => x"f8",
          2718 => x"11",
          2719 => x"82",
          2720 => x"f8",
          2721 => x"d6",
          2722 => x"05",
          2723 => x"89",
          2724 => x"80",
          2725 => x"e4",
          2726 => x"0c",
          2727 => x"82",
          2728 => x"f8",
          2729 => x"d6",
          2730 => x"05",
          2731 => x"72",
          2732 => x"38",
          2733 => x"d6",
          2734 => x"05",
          2735 => x"39",
          2736 => x"08",
          2737 => x"70",
          2738 => x"08",
          2739 => x"29",
          2740 => x"08",
          2741 => x"70",
          2742 => x"e4",
          2743 => x"0c",
          2744 => x"08",
          2745 => x"70",
          2746 => x"71",
          2747 => x"51",
          2748 => x"53",
          2749 => x"d6",
          2750 => x"05",
          2751 => x"39",
          2752 => x"08",
          2753 => x"53",
          2754 => x"90",
          2755 => x"e4",
          2756 => x"08",
          2757 => x"e4",
          2758 => x"0c",
          2759 => x"08",
          2760 => x"82",
          2761 => x"fc",
          2762 => x"0c",
          2763 => x"82",
          2764 => x"ec",
          2765 => x"d6",
          2766 => x"05",
          2767 => x"d8",
          2768 => x"0d",
          2769 => x"0c",
          2770 => x"0d",
          2771 => x"70",
          2772 => x"74",
          2773 => x"df",
          2774 => x"77",
          2775 => x"85",
          2776 => x"80",
          2777 => x"33",
          2778 => x"2e",
          2779 => x"86",
          2780 => x"55",
          2781 => x"57",
          2782 => x"82",
          2783 => x"70",
          2784 => x"e5",
          2785 => x"d6",
          2786 => x"d6",
          2787 => x"75",
          2788 => x"52",
          2789 => x"3f",
          2790 => x"08",
          2791 => x"16",
          2792 => x"81",
          2793 => x"38",
          2794 => x"81",
          2795 => x"54",
          2796 => x"c4",
          2797 => x"73",
          2798 => x"0c",
          2799 => x"04",
          2800 => x"73",
          2801 => x"26",
          2802 => x"71",
          2803 => x"ac",
          2804 => x"71",
          2805 => x"b2",
          2806 => x"80",
          2807 => x"d8",
          2808 => x"39",
          2809 => x"51",
          2810 => x"82",
          2811 => x"80",
          2812 => x"b3",
          2813 => x"e4",
          2814 => x"98",
          2815 => x"39",
          2816 => x"51",
          2817 => x"82",
          2818 => x"80",
          2819 => x"b3",
          2820 => x"c8",
          2821 => x"ec",
          2822 => x"39",
          2823 => x"51",
          2824 => x"b4",
          2825 => x"39",
          2826 => x"51",
          2827 => x"b4",
          2828 => x"39",
          2829 => x"51",
          2830 => x"b5",
          2831 => x"39",
          2832 => x"51",
          2833 => x"b5",
          2834 => x"39",
          2835 => x"51",
          2836 => x"b5",
          2837 => x"39",
          2838 => x"51",
          2839 => x"83",
          2840 => x"fb",
          2841 => x"79",
          2842 => x"87",
          2843 => x"38",
          2844 => x"87",
          2845 => x"90",
          2846 => x"52",
          2847 => x"af",
          2848 => x"d8",
          2849 => x"51",
          2850 => x"82",
          2851 => x"54",
          2852 => x"52",
          2853 => x"51",
          2854 => x"3f",
          2855 => x"04",
          2856 => x"66",
          2857 => x"80",
          2858 => x"5b",
          2859 => x"78",
          2860 => x"07",
          2861 => x"57",
          2862 => x"56",
          2863 => x"26",
          2864 => x"56",
          2865 => x"70",
          2866 => x"51",
          2867 => x"74",
          2868 => x"81",
          2869 => x"8c",
          2870 => x"56",
          2871 => x"3f",
          2872 => x"08",
          2873 => x"d8",
          2874 => x"82",
          2875 => x"87",
          2876 => x"0c",
          2877 => x"08",
          2878 => x"d4",
          2879 => x"80",
          2880 => x"75",
          2881 => x"8b",
          2882 => x"d8",
          2883 => x"d6",
          2884 => x"38",
          2885 => x"80",
          2886 => x"74",
          2887 => x"59",
          2888 => x"96",
          2889 => x"51",
          2890 => x"3f",
          2891 => x"78",
          2892 => x"7b",
          2893 => x"2a",
          2894 => x"57",
          2895 => x"80",
          2896 => x"82",
          2897 => x"87",
          2898 => x"08",
          2899 => x"fe",
          2900 => x"56",
          2901 => x"d8",
          2902 => x"0d",
          2903 => x"0d",
          2904 => x"05",
          2905 => x"59",
          2906 => x"80",
          2907 => x"7b",
          2908 => x"3f",
          2909 => x"08",
          2910 => x"77",
          2911 => x"38",
          2912 => x"bf",
          2913 => x"82",
          2914 => x"82",
          2915 => x"82",
          2916 => x"82",
          2917 => x"54",
          2918 => x"08",
          2919 => x"b8",
          2920 => x"b6",
          2921 => x"b8",
          2922 => x"f2",
          2923 => x"55",
          2924 => x"d6",
          2925 => x"52",
          2926 => x"2d",
          2927 => x"08",
          2928 => x"79",
          2929 => x"d6",
          2930 => x"3d",
          2931 => x"3d",
          2932 => x"63",
          2933 => x"80",
          2934 => x"73",
          2935 => x"41",
          2936 => x"5e",
          2937 => x"52",
          2938 => x"51",
          2939 => x"3f",
          2940 => x"51",
          2941 => x"3f",
          2942 => x"79",
          2943 => x"38",
          2944 => x"89",
          2945 => x"2e",
          2946 => x"c6",
          2947 => x"53",
          2948 => x"8e",
          2949 => x"52",
          2950 => x"51",
          2951 => x"3f",
          2952 => x"b6",
          2953 => x"b7",
          2954 => x"15",
          2955 => x"39",
          2956 => x"72",
          2957 => x"38",
          2958 => x"82",
          2959 => x"ff",
          2960 => x"89",
          2961 => x"f4",
          2962 => x"8d",
          2963 => x"55",
          2964 => x"18",
          2965 => x"27",
          2966 => x"33",
          2967 => x"80",
          2968 => x"f5",
          2969 => x"82",
          2970 => x"ff",
          2971 => x"81",
          2972 => x"f2",
          2973 => x"a0",
          2974 => x"3f",
          2975 => x"82",
          2976 => x"ff",
          2977 => x"80",
          2978 => x"27",
          2979 => x"74",
          2980 => x"55",
          2981 => x"72",
          2982 => x"38",
          2983 => x"53",
          2984 => x"83",
          2985 => x"75",
          2986 => x"81",
          2987 => x"53",
          2988 => x"90",
          2989 => x"fe",
          2990 => x"82",
          2991 => x"52",
          2992 => x"39",
          2993 => x"08",
          2994 => x"d5",
          2995 => x"15",
          2996 => x"39",
          2997 => x"51",
          2998 => x"78",
          2999 => x"5c",
          3000 => x"3f",
          3001 => x"08",
          3002 => x"98",
          3003 => x"76",
          3004 => x"81",
          3005 => x"9c",
          3006 => x"d6",
          3007 => x"2b",
          3008 => x"70",
          3009 => x"30",
          3010 => x"70",
          3011 => x"07",
          3012 => x"06",
          3013 => x"59",
          3014 => x"80",
          3015 => x"38",
          3016 => x"09",
          3017 => x"38",
          3018 => x"39",
          3019 => x"72",
          3020 => x"b2",
          3021 => x"72",
          3022 => x"0c",
          3023 => x"04",
          3024 => x"02",
          3025 => x"82",
          3026 => x"82",
          3027 => x"55",
          3028 => x"3f",
          3029 => x"22",
          3030 => x"3f",
          3031 => x"54",
          3032 => x"53",
          3033 => x"33",
          3034 => x"b8",
          3035 => x"e9",
          3036 => x"2e",
          3037 => x"f4",
          3038 => x"0d",
          3039 => x"0d",
          3040 => x"80",
          3041 => x"dc",
          3042 => x"99",
          3043 => x"b7",
          3044 => x"ce",
          3045 => x"99",
          3046 => x"81",
          3047 => x"06",
          3048 => x"80",
          3049 => x"81",
          3050 => x"3f",
          3051 => x"51",
          3052 => x"80",
          3053 => x"3f",
          3054 => x"70",
          3055 => x"52",
          3056 => x"92",
          3057 => x"99",
          3058 => x"b7",
          3059 => x"92",
          3060 => x"98",
          3061 => x"83",
          3062 => x"06",
          3063 => x"80",
          3064 => x"81",
          3065 => x"3f",
          3066 => x"51",
          3067 => x"80",
          3068 => x"3f",
          3069 => x"70",
          3070 => x"52",
          3071 => x"92",
          3072 => x"98",
          3073 => x"b8",
          3074 => x"d6",
          3075 => x"98",
          3076 => x"85",
          3077 => x"06",
          3078 => x"80",
          3079 => x"81",
          3080 => x"3f",
          3081 => x"51",
          3082 => x"80",
          3083 => x"3f",
          3084 => x"70",
          3085 => x"52",
          3086 => x"92",
          3087 => x"98",
          3088 => x"b8",
          3089 => x"9a",
          3090 => x"97",
          3091 => x"87",
          3092 => x"06",
          3093 => x"80",
          3094 => x"81",
          3095 => x"3f",
          3096 => x"51",
          3097 => x"80",
          3098 => x"3f",
          3099 => x"70",
          3100 => x"52",
          3101 => x"92",
          3102 => x"97",
          3103 => x"b8",
          3104 => x"de",
          3105 => x"97",
          3106 => x"e0",
          3107 => x"0d",
          3108 => x"0d",
          3109 => x"05",
          3110 => x"70",
          3111 => x"80",
          3112 => x"e2",
          3113 => x"0b",
          3114 => x"33",
          3115 => x"38",
          3116 => x"b9",
          3117 => x"ed",
          3118 => x"8a",
          3119 => x"d6",
          3120 => x"70",
          3121 => x"08",
          3122 => x"82",
          3123 => x"51",
          3124 => x"0b",
          3125 => x"34",
          3126 => x"d0",
          3127 => x"73",
          3128 => x"81",
          3129 => x"82",
          3130 => x"74",
          3131 => x"81",
          3132 => x"82",
          3133 => x"80",
          3134 => x"82",
          3135 => x"51",
          3136 => x"91",
          3137 => x"e8",
          3138 => x"a1",
          3139 => x"0b",
          3140 => x"c8",
          3141 => x"82",
          3142 => x"54",
          3143 => x"09",
          3144 => x"38",
          3145 => x"53",
          3146 => x"51",
          3147 => x"80",
          3148 => x"d8",
          3149 => x"0d",
          3150 => x"0d",
          3151 => x"5e",
          3152 => x"ed",
          3153 => x"81",
          3154 => x"80",
          3155 => x"82",
          3156 => x"81",
          3157 => x"78",
          3158 => x"81",
          3159 => x"97",
          3160 => x"53",
          3161 => x"52",
          3162 => x"fa",
          3163 => x"78",
          3164 => x"84",
          3165 => x"d5",
          3166 => x"d8",
          3167 => x"88",
          3168 => x"c8",
          3169 => x"39",
          3170 => x"5e",
          3171 => x"51",
          3172 => x"3f",
          3173 => x"47",
          3174 => x"52",
          3175 => x"f1",
          3176 => x"ff",
          3177 => x"f3",
          3178 => x"d6",
          3179 => x"2b",
          3180 => x"51",
          3181 => x"c2",
          3182 => x"38",
          3183 => x"24",
          3184 => x"bd",
          3185 => x"38",
          3186 => x"90",
          3187 => x"2e",
          3188 => x"78",
          3189 => x"da",
          3190 => x"39",
          3191 => x"2e",
          3192 => x"78",
          3193 => x"85",
          3194 => x"bf",
          3195 => x"38",
          3196 => x"78",
          3197 => x"89",
          3198 => x"80",
          3199 => x"38",
          3200 => x"2e",
          3201 => x"78",
          3202 => x"89",
          3203 => x"a1",
          3204 => x"83",
          3205 => x"38",
          3206 => x"24",
          3207 => x"81",
          3208 => x"ed",
          3209 => x"39",
          3210 => x"2e",
          3211 => x"8a",
          3212 => x"3d",
          3213 => x"53",
          3214 => x"51",
          3215 => x"82",
          3216 => x"80",
          3217 => x"38",
          3218 => x"fc",
          3219 => x"84",
          3220 => x"a4",
          3221 => x"d8",
          3222 => x"fe",
          3223 => x"3d",
          3224 => x"53",
          3225 => x"51",
          3226 => x"82",
          3227 => x"86",
          3228 => x"d8",
          3229 => x"ba",
          3230 => x"ae",
          3231 => x"64",
          3232 => x"7b",
          3233 => x"38",
          3234 => x"7a",
          3235 => x"5c",
          3236 => x"26",
          3237 => x"db",
          3238 => x"ff",
          3239 => x"ff",
          3240 => x"eb",
          3241 => x"d6",
          3242 => x"2e",
          3243 => x"b5",
          3244 => x"11",
          3245 => x"05",
          3246 => x"3f",
          3247 => x"08",
          3248 => x"c8",
          3249 => x"fe",
          3250 => x"ff",
          3251 => x"eb",
          3252 => x"d6",
          3253 => x"2e",
          3254 => x"82",
          3255 => x"ff",
          3256 => x"64",
          3257 => x"27",
          3258 => x"62",
          3259 => x"81",
          3260 => x"79",
          3261 => x"05",
          3262 => x"b5",
          3263 => x"11",
          3264 => x"05",
          3265 => x"3f",
          3266 => x"08",
          3267 => x"fc",
          3268 => x"fe",
          3269 => x"ff",
          3270 => x"ea",
          3271 => x"d6",
          3272 => x"2e",
          3273 => x"b5",
          3274 => x"11",
          3275 => x"05",
          3276 => x"3f",
          3277 => x"08",
          3278 => x"d0",
          3279 => x"a0",
          3280 => x"95",
          3281 => x"79",
          3282 => x"38",
          3283 => x"7b",
          3284 => x"5b",
          3285 => x"92",
          3286 => x"7a",
          3287 => x"53",
          3288 => x"ba",
          3289 => x"ac",
          3290 => x"1a",
          3291 => x"44",
          3292 => x"8a",
          3293 => x"3f",
          3294 => x"b5",
          3295 => x"11",
          3296 => x"05",
          3297 => x"3f",
          3298 => x"08",
          3299 => x"82",
          3300 => x"59",
          3301 => x"89",
          3302 => x"f0",
          3303 => x"cd",
          3304 => x"b9",
          3305 => x"80",
          3306 => x"82",
          3307 => x"45",
          3308 => x"d4",
          3309 => x"78",
          3310 => x"38",
          3311 => x"08",
          3312 => x"82",
          3313 => x"59",
          3314 => x"88",
          3315 => x"88",
          3316 => x"39",
          3317 => x"33",
          3318 => x"2e",
          3319 => x"d4",
          3320 => x"89",
          3321 => x"a0",
          3322 => x"05",
          3323 => x"fe",
          3324 => x"ff",
          3325 => x"e8",
          3326 => x"d6",
          3327 => x"de",
          3328 => x"b8",
          3329 => x"80",
          3330 => x"82",
          3331 => x"44",
          3332 => x"82",
          3333 => x"59",
          3334 => x"88",
          3335 => x"fc",
          3336 => x"39",
          3337 => x"33",
          3338 => x"2e",
          3339 => x"d4",
          3340 => x"aa",
          3341 => x"bb",
          3342 => x"80",
          3343 => x"82",
          3344 => x"44",
          3345 => x"d4",
          3346 => x"78",
          3347 => x"38",
          3348 => x"08",
          3349 => x"82",
          3350 => x"88",
          3351 => x"3d",
          3352 => x"53",
          3353 => x"51",
          3354 => x"82",
          3355 => x"80",
          3356 => x"80",
          3357 => x"7a",
          3358 => x"38",
          3359 => x"90",
          3360 => x"70",
          3361 => x"2a",
          3362 => x"51",
          3363 => x"78",
          3364 => x"38",
          3365 => x"83",
          3366 => x"82",
          3367 => x"c6",
          3368 => x"55",
          3369 => x"53",
          3370 => x"51",
          3371 => x"82",
          3372 => x"87",
          3373 => x"3d",
          3374 => x"53",
          3375 => x"51",
          3376 => x"82",
          3377 => x"80",
          3378 => x"38",
          3379 => x"fc",
          3380 => x"84",
          3381 => x"a0",
          3382 => x"d8",
          3383 => x"a4",
          3384 => x"02",
          3385 => x"33",
          3386 => x"81",
          3387 => x"3d",
          3388 => x"53",
          3389 => x"51",
          3390 => x"82",
          3391 => x"e1",
          3392 => x"39",
          3393 => x"54",
          3394 => x"e4",
          3395 => x"c9",
          3396 => x"b8",
          3397 => x"f8",
          3398 => x"ff",
          3399 => x"79",
          3400 => x"59",
          3401 => x"f8",
          3402 => x"79",
          3403 => x"b5",
          3404 => x"11",
          3405 => x"05",
          3406 => x"3f",
          3407 => x"08",
          3408 => x"38",
          3409 => x"80",
          3410 => x"79",
          3411 => x"05",
          3412 => x"39",
          3413 => x"51",
          3414 => x"ff",
          3415 => x"3d",
          3416 => x"53",
          3417 => x"51",
          3418 => x"82",
          3419 => x"80",
          3420 => x"38",
          3421 => x"f0",
          3422 => x"84",
          3423 => x"a7",
          3424 => x"d8",
          3425 => x"a6",
          3426 => x"02",
          3427 => x"22",
          3428 => x"05",
          3429 => x"42",
          3430 => x"f0",
          3431 => x"84",
          3432 => x"83",
          3433 => x"d8",
          3434 => x"f7",
          3435 => x"70",
          3436 => x"82",
          3437 => x"ff",
          3438 => x"82",
          3439 => x"53",
          3440 => x"79",
          3441 => x"e6",
          3442 => x"79",
          3443 => x"ae",
          3444 => x"38",
          3445 => x"87",
          3446 => x"05",
          3447 => x"b5",
          3448 => x"11",
          3449 => x"05",
          3450 => x"3f",
          3451 => x"08",
          3452 => x"38",
          3453 => x"80",
          3454 => x"79",
          3455 => x"5b",
          3456 => x"ff",
          3457 => x"ba",
          3458 => x"d8",
          3459 => x"39",
          3460 => x"f4",
          3461 => x"84",
          3462 => x"8b",
          3463 => x"d8",
          3464 => x"f6",
          3465 => x"3d",
          3466 => x"53",
          3467 => x"51",
          3468 => x"82",
          3469 => x"80",
          3470 => x"61",
          3471 => x"59",
          3472 => x"42",
          3473 => x"f0",
          3474 => x"84",
          3475 => x"d7",
          3476 => x"d8",
          3477 => x"f6",
          3478 => x"70",
          3479 => x"82",
          3480 => x"ff",
          3481 => x"82",
          3482 => x"53",
          3483 => x"79",
          3484 => x"ba",
          3485 => x"79",
          3486 => x"ae",
          3487 => x"38",
          3488 => x"9b",
          3489 => x"fe",
          3490 => x"ff",
          3491 => x"de",
          3492 => x"d6",
          3493 => x"2e",
          3494 => x"61",
          3495 => x"61",
          3496 => x"ff",
          3497 => x"ba",
          3498 => x"b8",
          3499 => x"39",
          3500 => x"80",
          3501 => x"84",
          3502 => x"bc",
          3503 => x"d8",
          3504 => x"f5",
          3505 => x"52",
          3506 => x"51",
          3507 => x"3f",
          3508 => x"04",
          3509 => x"80",
          3510 => x"84",
          3511 => x"98",
          3512 => x"d8",
          3513 => x"f5",
          3514 => x"52",
          3515 => x"51",
          3516 => x"3f",
          3517 => x"2d",
          3518 => x"08",
          3519 => x"8c",
          3520 => x"d8",
          3521 => x"bb",
          3522 => x"a5",
          3523 => x"fc",
          3524 => x"e4",
          3525 => x"3f",
          3526 => x"3f",
          3527 => x"82",
          3528 => x"c1",
          3529 => x"59",
          3530 => x"91",
          3531 => x"dc",
          3532 => x"33",
          3533 => x"2e",
          3534 => x"80",
          3535 => x"51",
          3536 => x"82",
          3537 => x"5d",
          3538 => x"08",
          3539 => x"92",
          3540 => x"d8",
          3541 => x"3d",
          3542 => x"51",
          3543 => x"82",
          3544 => x"60",
          3545 => x"5c",
          3546 => x"81",
          3547 => x"d6",
          3548 => x"cd",
          3549 => x"d6",
          3550 => x"26",
          3551 => x"81",
          3552 => x"2e",
          3553 => x"82",
          3554 => x"7a",
          3555 => x"38",
          3556 => x"7a",
          3557 => x"38",
          3558 => x"82",
          3559 => x"7b",
          3560 => x"98",
          3561 => x"82",
          3562 => x"b5",
          3563 => x"05",
          3564 => x"8d",
          3565 => x"7b",
          3566 => x"ff",
          3567 => x"cd",
          3568 => x"39",
          3569 => x"bc",
          3570 => x"53",
          3571 => x"52",
          3572 => x"b0",
          3573 => x"a6",
          3574 => x"39",
          3575 => x"53",
          3576 => x"52",
          3577 => x"b0",
          3578 => x"a6",
          3579 => x"d3",
          3580 => x"d7",
          3581 => x"56",
          3582 => x"54",
          3583 => x"53",
          3584 => x"52",
          3585 => x"b0",
          3586 => x"d1",
          3587 => x"d8",
          3588 => x"d8",
          3589 => x"30",
          3590 => x"80",
          3591 => x"5b",
          3592 => x"7a",
          3593 => x"38",
          3594 => x"7a",
          3595 => x"80",
          3596 => x"81",
          3597 => x"ff",
          3598 => x"7a",
          3599 => x"7f",
          3600 => x"81",
          3601 => x"78",
          3602 => x"ff",
          3603 => x"06",
          3604 => x"bc",
          3605 => x"bf",
          3606 => x"51",
          3607 => x"f2",
          3608 => x"bc",
          3609 => x"be",
          3610 => x"a0",
          3611 => x"0d",
          3612 => x"d7",
          3613 => x"c0",
          3614 => x"53",
          3615 => x"52",
          3616 => x"ab",
          3617 => x"d8",
          3618 => x"87",
          3619 => x"08",
          3620 => x"84",
          3621 => x"51",
          3622 => x"72",
          3623 => x"08",
          3624 => x"94",
          3625 => x"c0",
          3626 => x"53",
          3627 => x"52",
          3628 => x"fb",
          3629 => x"d8",
          3630 => x"87",
          3631 => x"08",
          3632 => x"84",
          3633 => x"51",
          3634 => x"72",
          3635 => x"08",
          3636 => x"94",
          3637 => x"80",
          3638 => x"c0",
          3639 => x"8c",
          3640 => x"87",
          3641 => x"0c",
          3642 => x"80",
          3643 => x"70",
          3644 => x"0c",
          3645 => x"fe",
          3646 => x"38",
          3647 => x"80",
          3648 => x"c5",
          3649 => x"70",
          3650 => x"0c",
          3651 => x"fe",
          3652 => x"38",
          3653 => x"c8",
          3654 => x"3f",
          3655 => x"c5",
          3656 => x"3f",
          3657 => x"cc",
          3658 => x"3f",
          3659 => x"cc",
          3660 => x"3f",
          3661 => x"cf",
          3662 => x"3f",
          3663 => x"51",
          3664 => x"80",
          3665 => x"a6",
          3666 => x"99",
          3667 => x"9a",
          3668 => x"02",
          3669 => x"05",
          3670 => x"85",
          3671 => x"f2",
          3672 => x"82",
          3673 => x"82",
          3674 => x"82",
          3675 => x"ff",
          3676 => x"88",
          3677 => x"ec",
          3678 => x"8c",
          3679 => x"e4",
          3680 => x"98",
          3681 => x"dc",
          3682 => x"fc",
          3683 => x"3f",
          3684 => x"ac",
          3685 => x"3f",
          3686 => x"3d",
          3687 => x"83",
          3688 => x"2b",
          3689 => x"3f",
          3690 => x"08",
          3691 => x"72",
          3692 => x"54",
          3693 => x"25",
          3694 => x"82",
          3695 => x"84",
          3696 => x"fc",
          3697 => x"70",
          3698 => x"80",
          3699 => x"72",
          3700 => x"8a",
          3701 => x"51",
          3702 => x"09",
          3703 => x"38",
          3704 => x"f1",
          3705 => x"51",
          3706 => x"09",
          3707 => x"38",
          3708 => x"81",
          3709 => x"73",
          3710 => x"81",
          3711 => x"84",
          3712 => x"52",
          3713 => x"52",
          3714 => x"2e",
          3715 => x"54",
          3716 => x"9d",
          3717 => x"38",
          3718 => x"12",
          3719 => x"33",
          3720 => x"a0",
          3721 => x"81",
          3722 => x"2e",
          3723 => x"ea",
          3724 => x"33",
          3725 => x"a0",
          3726 => x"06",
          3727 => x"54",
          3728 => x"70",
          3729 => x"25",
          3730 => x"51",
          3731 => x"2e",
          3732 => x"72",
          3733 => x"54",
          3734 => x"0c",
          3735 => x"82",
          3736 => x"86",
          3737 => x"fc",
          3738 => x"53",
          3739 => x"2e",
          3740 => x"3d",
          3741 => x"72",
          3742 => x"3f",
          3743 => x"08",
          3744 => x"53",
          3745 => x"53",
          3746 => x"d8",
          3747 => x"0d",
          3748 => x"0d",
          3749 => x"33",
          3750 => x"53",
          3751 => x"8b",
          3752 => x"38",
          3753 => x"ff",
          3754 => x"52",
          3755 => x"81",
          3756 => x"13",
          3757 => x"52",
          3758 => x"80",
          3759 => x"13",
          3760 => x"52",
          3761 => x"80",
          3762 => x"13",
          3763 => x"52",
          3764 => x"80",
          3765 => x"13",
          3766 => x"52",
          3767 => x"26",
          3768 => x"8a",
          3769 => x"87",
          3770 => x"e7",
          3771 => x"38",
          3772 => x"c0",
          3773 => x"72",
          3774 => x"98",
          3775 => x"13",
          3776 => x"98",
          3777 => x"13",
          3778 => x"98",
          3779 => x"13",
          3780 => x"98",
          3781 => x"13",
          3782 => x"98",
          3783 => x"13",
          3784 => x"98",
          3785 => x"87",
          3786 => x"0c",
          3787 => x"98",
          3788 => x"0b",
          3789 => x"9c",
          3790 => x"71",
          3791 => x"0c",
          3792 => x"04",
          3793 => x"7f",
          3794 => x"98",
          3795 => x"7d",
          3796 => x"98",
          3797 => x"7d",
          3798 => x"c0",
          3799 => x"5a",
          3800 => x"34",
          3801 => x"b4",
          3802 => x"83",
          3803 => x"c0",
          3804 => x"5a",
          3805 => x"34",
          3806 => x"ac",
          3807 => x"85",
          3808 => x"c0",
          3809 => x"5a",
          3810 => x"34",
          3811 => x"a4",
          3812 => x"88",
          3813 => x"c0",
          3814 => x"5a",
          3815 => x"23",
          3816 => x"79",
          3817 => x"06",
          3818 => x"ff",
          3819 => x"86",
          3820 => x"85",
          3821 => x"84",
          3822 => x"83",
          3823 => x"82",
          3824 => x"7d",
          3825 => x"06",
          3826 => x"b0",
          3827 => x"89",
          3828 => x"0d",
          3829 => x"0d",
          3830 => x"33",
          3831 => x"33",
          3832 => x"06",
          3833 => x"87",
          3834 => x"51",
          3835 => x"86",
          3836 => x"94",
          3837 => x"08",
          3838 => x"70",
          3839 => x"54",
          3840 => x"2e",
          3841 => x"91",
          3842 => x"06",
          3843 => x"d7",
          3844 => x"32",
          3845 => x"51",
          3846 => x"2e",
          3847 => x"93",
          3848 => x"06",
          3849 => x"ff",
          3850 => x"81",
          3851 => x"87",
          3852 => x"52",
          3853 => x"86",
          3854 => x"94",
          3855 => x"72",
          3856 => x"d6",
          3857 => x"3d",
          3858 => x"3d",
          3859 => x"05",
          3860 => x"70",
          3861 => x"52",
          3862 => x"d3",
          3863 => x"3d",
          3864 => x"3d",
          3865 => x"80",
          3866 => x"81",
          3867 => x"53",
          3868 => x"2e",
          3869 => x"71",
          3870 => x"81",
          3871 => x"ec",
          3872 => x"ff",
          3873 => x"55",
          3874 => x"94",
          3875 => x"80",
          3876 => x"87",
          3877 => x"51",
          3878 => x"96",
          3879 => x"06",
          3880 => x"70",
          3881 => x"38",
          3882 => x"70",
          3883 => x"51",
          3884 => x"72",
          3885 => x"81",
          3886 => x"70",
          3887 => x"38",
          3888 => x"70",
          3889 => x"51",
          3890 => x"38",
          3891 => x"06",
          3892 => x"94",
          3893 => x"80",
          3894 => x"87",
          3895 => x"52",
          3896 => x"81",
          3897 => x"70",
          3898 => x"53",
          3899 => x"ff",
          3900 => x"82",
          3901 => x"89",
          3902 => x"fe",
          3903 => x"d3",
          3904 => x"81",
          3905 => x"52",
          3906 => x"84",
          3907 => x"2e",
          3908 => x"c0",
          3909 => x"70",
          3910 => x"2a",
          3911 => x"51",
          3912 => x"80",
          3913 => x"71",
          3914 => x"51",
          3915 => x"80",
          3916 => x"2e",
          3917 => x"c0",
          3918 => x"71",
          3919 => x"ff",
          3920 => x"d8",
          3921 => x"3d",
          3922 => x"3d",
          3923 => x"ec",
          3924 => x"ff",
          3925 => x"87",
          3926 => x"52",
          3927 => x"86",
          3928 => x"94",
          3929 => x"08",
          3930 => x"70",
          3931 => x"51",
          3932 => x"70",
          3933 => x"38",
          3934 => x"06",
          3935 => x"94",
          3936 => x"80",
          3937 => x"87",
          3938 => x"52",
          3939 => x"98",
          3940 => x"2c",
          3941 => x"71",
          3942 => x"0c",
          3943 => x"04",
          3944 => x"87",
          3945 => x"08",
          3946 => x"8a",
          3947 => x"70",
          3948 => x"b4",
          3949 => x"9e",
          3950 => x"d3",
          3951 => x"c0",
          3952 => x"82",
          3953 => x"87",
          3954 => x"08",
          3955 => x"0c",
          3956 => x"98",
          3957 => x"fc",
          3958 => x"9e",
          3959 => x"d4",
          3960 => x"c0",
          3961 => x"82",
          3962 => x"87",
          3963 => x"08",
          3964 => x"0c",
          3965 => x"b0",
          3966 => x"8c",
          3967 => x"9e",
          3968 => x"d4",
          3969 => x"c0",
          3970 => x"82",
          3971 => x"87",
          3972 => x"08",
          3973 => x"0c",
          3974 => x"c0",
          3975 => x"9c",
          3976 => x"9e",
          3977 => x"d4",
          3978 => x"c0",
          3979 => x"51",
          3980 => x"a4",
          3981 => x"9e",
          3982 => x"d4",
          3983 => x"c0",
          3984 => x"82",
          3985 => x"87",
          3986 => x"08",
          3987 => x"0c",
          3988 => x"d4",
          3989 => x"0b",
          3990 => x"90",
          3991 => x"80",
          3992 => x"52",
          3993 => x"2e",
          3994 => x"52",
          3995 => x"b5",
          3996 => x"87",
          3997 => x"08",
          3998 => x"0a",
          3999 => x"52",
          4000 => x"83",
          4001 => x"71",
          4002 => x"34",
          4003 => x"c0",
          4004 => x"70",
          4005 => x"06",
          4006 => x"70",
          4007 => x"38",
          4008 => x"82",
          4009 => x"80",
          4010 => x"9e",
          4011 => x"88",
          4012 => x"51",
          4013 => x"80",
          4014 => x"81",
          4015 => x"d4",
          4016 => x"0b",
          4017 => x"90",
          4018 => x"80",
          4019 => x"52",
          4020 => x"2e",
          4021 => x"52",
          4022 => x"b9",
          4023 => x"87",
          4024 => x"08",
          4025 => x"80",
          4026 => x"52",
          4027 => x"83",
          4028 => x"71",
          4029 => x"34",
          4030 => x"c0",
          4031 => x"70",
          4032 => x"06",
          4033 => x"70",
          4034 => x"38",
          4035 => x"82",
          4036 => x"80",
          4037 => x"9e",
          4038 => x"82",
          4039 => x"51",
          4040 => x"80",
          4041 => x"81",
          4042 => x"d4",
          4043 => x"0b",
          4044 => x"90",
          4045 => x"80",
          4046 => x"52",
          4047 => x"2e",
          4048 => x"52",
          4049 => x"bd",
          4050 => x"87",
          4051 => x"08",
          4052 => x"80",
          4053 => x"52",
          4054 => x"83",
          4055 => x"71",
          4056 => x"34",
          4057 => x"c0",
          4058 => x"70",
          4059 => x"51",
          4060 => x"80",
          4061 => x"81",
          4062 => x"d4",
          4063 => x"c0",
          4064 => x"70",
          4065 => x"70",
          4066 => x"51",
          4067 => x"d4",
          4068 => x"0b",
          4069 => x"90",
          4070 => x"80",
          4071 => x"52",
          4072 => x"83",
          4073 => x"71",
          4074 => x"34",
          4075 => x"90",
          4076 => x"f0",
          4077 => x"2a",
          4078 => x"70",
          4079 => x"34",
          4080 => x"c0",
          4081 => x"70",
          4082 => x"52",
          4083 => x"2e",
          4084 => x"52",
          4085 => x"c3",
          4086 => x"9e",
          4087 => x"87",
          4088 => x"70",
          4089 => x"34",
          4090 => x"04",
          4091 => x"82",
          4092 => x"ff",
          4093 => x"82",
          4094 => x"54",
          4095 => x"89",
          4096 => x"dc",
          4097 => x"d1",
          4098 => x"f0",
          4099 => x"d4",
          4100 => x"b6",
          4101 => x"80",
          4102 => x"82",
          4103 => x"82",
          4104 => x"11",
          4105 => x"be",
          4106 => x"93",
          4107 => x"d4",
          4108 => x"73",
          4109 => x"38",
          4110 => x"08",
          4111 => x"08",
          4112 => x"82",
          4113 => x"ff",
          4114 => x"82",
          4115 => x"54",
          4116 => x"94",
          4117 => x"f0",
          4118 => x"f4",
          4119 => x"52",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"33",
          4123 => x"2e",
          4124 => x"d3",
          4125 => x"d3",
          4126 => x"54",
          4127 => x"dc",
          4128 => x"d5",
          4129 => x"ba",
          4130 => x"80",
          4131 => x"82",
          4132 => x"82",
          4133 => x"11",
          4134 => x"be",
          4135 => x"92",
          4136 => x"d4",
          4137 => x"73",
          4138 => x"38",
          4139 => x"33",
          4140 => x"94",
          4141 => x"a1",
          4142 => x"c3",
          4143 => x"80",
          4144 => x"82",
          4145 => x"52",
          4146 => x"51",
          4147 => x"3f",
          4148 => x"33",
          4149 => x"2e",
          4150 => x"d4",
          4151 => x"82",
          4152 => x"ff",
          4153 => x"82",
          4154 => x"54",
          4155 => x"89",
          4156 => x"f4",
          4157 => x"ec",
          4158 => x"b7",
          4159 => x"80",
          4160 => x"82",
          4161 => x"ff",
          4162 => x"82",
          4163 => x"54",
          4164 => x"89",
          4165 => x"94",
          4166 => x"c8",
          4167 => x"bd",
          4168 => x"80",
          4169 => x"82",
          4170 => x"ff",
          4171 => x"82",
          4172 => x"54",
          4173 => x"89",
          4174 => x"a8",
          4175 => x"a4",
          4176 => x"b0",
          4177 => x"9c",
          4178 => x"98",
          4179 => x"c0",
          4180 => x"91",
          4181 => x"d4",
          4182 => x"82",
          4183 => x"ff",
          4184 => x"82",
          4185 => x"52",
          4186 => x"51",
          4187 => x"3f",
          4188 => x"51",
          4189 => x"3f",
          4190 => x"22",
          4191 => x"bc",
          4192 => x"d5",
          4193 => x"a8",
          4194 => x"84",
          4195 => x"51",
          4196 => x"82",
          4197 => x"bd",
          4198 => x"76",
          4199 => x"54",
          4200 => x"08",
          4201 => x"e4",
          4202 => x"ad",
          4203 => x"bb",
          4204 => x"80",
          4205 => x"82",
          4206 => x"56",
          4207 => x"52",
          4208 => x"eb",
          4209 => x"d8",
          4210 => x"c0",
          4211 => x"31",
          4212 => x"d6",
          4213 => x"82",
          4214 => x"ff",
          4215 => x"82",
          4216 => x"54",
          4217 => x"a9",
          4218 => x"b0",
          4219 => x"84",
          4220 => x"51",
          4221 => x"82",
          4222 => x"bd",
          4223 => x"76",
          4224 => x"54",
          4225 => x"08",
          4226 => x"bc",
          4227 => x"c9",
          4228 => x"ff",
          4229 => x"87",
          4230 => x"fe",
          4231 => x"92",
          4232 => x"05",
          4233 => x"26",
          4234 => x"84",
          4235 => x"ac",
          4236 => x"08",
          4237 => x"e8",
          4238 => x"82",
          4239 => x"97",
          4240 => x"f8",
          4241 => x"82",
          4242 => x"8b",
          4243 => x"84",
          4244 => x"82",
          4245 => x"ff",
          4246 => x"84",
          4247 => x"71",
          4248 => x"04",
          4249 => x"c0",
          4250 => x"04",
          4251 => x"08",
          4252 => x"84",
          4253 => x"3d",
          4254 => x"2b",
          4255 => x"79",
          4256 => x"98",
          4257 => x"13",
          4258 => x"51",
          4259 => x"51",
          4260 => x"82",
          4261 => x"33",
          4262 => x"74",
          4263 => x"82",
          4264 => x"08",
          4265 => x"05",
          4266 => x"71",
          4267 => x"52",
          4268 => x"09",
          4269 => x"38",
          4270 => x"82",
          4271 => x"85",
          4272 => x"fb",
          4273 => x"02",
          4274 => x"05",
          4275 => x"55",
          4276 => x"80",
          4277 => x"82",
          4278 => x"52",
          4279 => x"ad",
          4280 => x"f2",
          4281 => x"a0",
          4282 => x"c7",
          4283 => x"bc",
          4284 => x"51",
          4285 => x"3f",
          4286 => x"05",
          4287 => x"34",
          4288 => x"06",
          4289 => x"77",
          4290 => x"cd",
          4291 => x"34",
          4292 => x"04",
          4293 => x"7c",
          4294 => x"b7",
          4295 => x"88",
          4296 => x"33",
          4297 => x"33",
          4298 => x"82",
          4299 => x"70",
          4300 => x"59",
          4301 => x"74",
          4302 => x"38",
          4303 => x"93",
          4304 => x"a4",
          4305 => x"29",
          4306 => x"05",
          4307 => x"54",
          4308 => x"9f",
          4309 => x"d6",
          4310 => x"0c",
          4311 => x"33",
          4312 => x"82",
          4313 => x"70",
          4314 => x"5a",
          4315 => x"a7",
          4316 => x"78",
          4317 => x"ff",
          4318 => x"82",
          4319 => x"81",
          4320 => x"82",
          4321 => x"74",
          4322 => x"55",
          4323 => x"87",
          4324 => x"82",
          4325 => x"77",
          4326 => x"38",
          4327 => x"08",
          4328 => x"2e",
          4329 => x"d5",
          4330 => x"74",
          4331 => x"3d",
          4332 => x"76",
          4333 => x"75",
          4334 => x"d7",
          4335 => x"a0",
          4336 => x"51",
          4337 => x"3f",
          4338 => x"08",
          4339 => x"ba",
          4340 => x"0d",
          4341 => x"0d",
          4342 => x"53",
          4343 => x"08",
          4344 => x"2e",
          4345 => x"51",
          4346 => x"80",
          4347 => x"14",
          4348 => x"54",
          4349 => x"e6",
          4350 => x"82",
          4351 => x"82",
          4352 => x"52",
          4353 => x"95",
          4354 => x"80",
          4355 => x"82",
          4356 => x"51",
          4357 => x"80",
          4358 => x"a0",
          4359 => x"0d",
          4360 => x"0d",
          4361 => x"52",
          4362 => x"08",
          4363 => x"bb",
          4364 => x"d8",
          4365 => x"38",
          4366 => x"08",
          4367 => x"52",
          4368 => x"52",
          4369 => x"eb",
          4370 => x"d8",
          4371 => x"ba",
          4372 => x"ff",
          4373 => x"82",
          4374 => x"55",
          4375 => x"d6",
          4376 => x"9d",
          4377 => x"d8",
          4378 => x"70",
          4379 => x"80",
          4380 => x"53",
          4381 => x"17",
          4382 => x"52",
          4383 => x"d9",
          4384 => x"2e",
          4385 => x"ff",
          4386 => x"3d",
          4387 => x"3d",
          4388 => x"08",
          4389 => x"5a",
          4390 => x"58",
          4391 => x"82",
          4392 => x"51",
          4393 => x"3f",
          4394 => x"08",
          4395 => x"ff",
          4396 => x"a0",
          4397 => x"80",
          4398 => x"3d",
          4399 => x"81",
          4400 => x"82",
          4401 => x"80",
          4402 => x"75",
          4403 => x"b6",
          4404 => x"d8",
          4405 => x"58",
          4406 => x"82",
          4407 => x"25",
          4408 => x"d6",
          4409 => x"05",
          4410 => x"55",
          4411 => x"74",
          4412 => x"70",
          4413 => x"2a",
          4414 => x"78",
          4415 => x"38",
          4416 => x"38",
          4417 => x"08",
          4418 => x"53",
          4419 => x"db",
          4420 => x"d8",
          4421 => x"89",
          4422 => x"94",
          4423 => x"b9",
          4424 => x"2e",
          4425 => x"9b",
          4426 => x"79",
          4427 => x"c4",
          4428 => x"ff",
          4429 => x"ab",
          4430 => x"82",
          4431 => x"74",
          4432 => x"77",
          4433 => x"0c",
          4434 => x"04",
          4435 => x"7c",
          4436 => x"71",
          4437 => x"59",
          4438 => x"a0",
          4439 => x"06",
          4440 => x"33",
          4441 => x"77",
          4442 => x"38",
          4443 => x"5b",
          4444 => x"56",
          4445 => x"a0",
          4446 => x"06",
          4447 => x"75",
          4448 => x"80",
          4449 => x"29",
          4450 => x"05",
          4451 => x"55",
          4452 => x"3f",
          4453 => x"08",
          4454 => x"74",
          4455 => x"b3",
          4456 => x"d6",
          4457 => x"c5",
          4458 => x"33",
          4459 => x"2e",
          4460 => x"82",
          4461 => x"b5",
          4462 => x"3f",
          4463 => x"1a",
          4464 => x"fc",
          4465 => x"05",
          4466 => x"3f",
          4467 => x"08",
          4468 => x"38",
          4469 => x"78",
          4470 => x"fd",
          4471 => x"d6",
          4472 => x"ff",
          4473 => x"85",
          4474 => x"91",
          4475 => x"70",
          4476 => x"51",
          4477 => x"27",
          4478 => x"80",
          4479 => x"d6",
          4480 => x"3d",
          4481 => x"3d",
          4482 => x"08",
          4483 => x"b4",
          4484 => x"5f",
          4485 => x"af",
          4486 => x"d5",
          4487 => x"d5",
          4488 => x"5b",
          4489 => x"38",
          4490 => x"9c",
          4491 => x"73",
          4492 => x"55",
          4493 => x"81",
          4494 => x"70",
          4495 => x"56",
          4496 => x"81",
          4497 => x"51",
          4498 => x"82",
          4499 => x"82",
          4500 => x"82",
          4501 => x"80",
          4502 => x"38",
          4503 => x"52",
          4504 => x"08",
          4505 => x"c6",
          4506 => x"d8",
          4507 => x"8c",
          4508 => x"c0",
          4509 => x"ec",
          4510 => x"39",
          4511 => x"08",
          4512 => x"a0",
          4513 => x"f8",
          4514 => x"70",
          4515 => x"9a",
          4516 => x"d6",
          4517 => x"82",
          4518 => x"74",
          4519 => x"06",
          4520 => x"82",
          4521 => x"51",
          4522 => x"3f",
          4523 => x"08",
          4524 => x"82",
          4525 => x"25",
          4526 => x"d6",
          4527 => x"05",
          4528 => x"55",
          4529 => x"80",
          4530 => x"ff",
          4531 => x"51",
          4532 => x"81",
          4533 => x"ff",
          4534 => x"93",
          4535 => x"38",
          4536 => x"ff",
          4537 => x"06",
          4538 => x"86",
          4539 => x"d5",
          4540 => x"8c",
          4541 => x"a0",
          4542 => x"84",
          4543 => x"3f",
          4544 => x"ec",
          4545 => x"d6",
          4546 => x"2b",
          4547 => x"51",
          4548 => x"2e",
          4549 => x"81",
          4550 => x"ee",
          4551 => x"98",
          4552 => x"2c",
          4553 => x"33",
          4554 => x"70",
          4555 => x"98",
          4556 => x"84",
          4557 => x"94",
          4558 => x"15",
          4559 => x"51",
          4560 => x"59",
          4561 => x"58",
          4562 => x"78",
          4563 => x"38",
          4564 => x"b4",
          4565 => x"80",
          4566 => x"ff",
          4567 => x"98",
          4568 => x"80",
          4569 => x"ce",
          4570 => x"74",
          4571 => x"f6",
          4572 => x"d6",
          4573 => x"ff",
          4574 => x"80",
          4575 => x"74",
          4576 => x"34",
          4577 => x"39",
          4578 => x"0a",
          4579 => x"0a",
          4580 => x"2c",
          4581 => x"06",
          4582 => x"73",
          4583 => x"38",
          4584 => x"52",
          4585 => x"ce",
          4586 => x"d8",
          4587 => x"06",
          4588 => x"38",
          4589 => x"56",
          4590 => x"80",
          4591 => x"1c",
          4592 => x"ee",
          4593 => x"98",
          4594 => x"2c",
          4595 => x"33",
          4596 => x"70",
          4597 => x"10",
          4598 => x"2b",
          4599 => x"11",
          4600 => x"51",
          4601 => x"51",
          4602 => x"2e",
          4603 => x"fe",
          4604 => x"c3",
          4605 => x"7d",
          4606 => x"82",
          4607 => x"80",
          4608 => x"90",
          4609 => x"75",
          4610 => x"34",
          4611 => x"90",
          4612 => x"3d",
          4613 => x"0c",
          4614 => x"95",
          4615 => x"38",
          4616 => x"82",
          4617 => x"54",
          4618 => x"82",
          4619 => x"54",
          4620 => x"fd",
          4621 => x"ee",
          4622 => x"73",
          4623 => x"38",
          4624 => x"70",
          4625 => x"55",
          4626 => x"9e",
          4627 => x"54",
          4628 => x"15",
          4629 => x"80",
          4630 => x"ff",
          4631 => x"98",
          4632 => x"9c",
          4633 => x"55",
          4634 => x"ee",
          4635 => x"11",
          4636 => x"82",
          4637 => x"73",
          4638 => x"3d",
          4639 => x"82",
          4640 => x"54",
          4641 => x"89",
          4642 => x"54",
          4643 => x"98",
          4644 => x"9c",
          4645 => x"80",
          4646 => x"ff",
          4647 => x"98",
          4648 => x"98",
          4649 => x"56",
          4650 => x"25",
          4651 => x"f2",
          4652 => x"74",
          4653 => x"52",
          4654 => x"f7",
          4655 => x"80",
          4656 => x"80",
          4657 => x"98",
          4658 => x"98",
          4659 => x"55",
          4660 => x"da",
          4661 => x"9c",
          4662 => x"2b",
          4663 => x"82",
          4664 => x"5a",
          4665 => x"74",
          4666 => x"94",
          4667 => x"bc",
          4668 => x"51",
          4669 => x"3f",
          4670 => x"0a",
          4671 => x"0a",
          4672 => x"2c",
          4673 => x"33",
          4674 => x"73",
          4675 => x"38",
          4676 => x"83",
          4677 => x"0b",
          4678 => x"82",
          4679 => x"80",
          4680 => x"a0",
          4681 => x"3f",
          4682 => x"82",
          4683 => x"70",
          4684 => x"55",
          4685 => x"2e",
          4686 => x"82",
          4687 => x"ff",
          4688 => x"82",
          4689 => x"ff",
          4690 => x"82",
          4691 => x"82",
          4692 => x"52",
          4693 => x"a0",
          4694 => x"ee",
          4695 => x"98",
          4696 => x"2c",
          4697 => x"33",
          4698 => x"57",
          4699 => x"ad",
          4700 => x"54",
          4701 => x"74",
          4702 => x"bc",
          4703 => x"33",
          4704 => x"af",
          4705 => x"80",
          4706 => x"80",
          4707 => x"98",
          4708 => x"98",
          4709 => x"55",
          4710 => x"d5",
          4711 => x"bc",
          4712 => x"51",
          4713 => x"3f",
          4714 => x"33",
          4715 => x"70",
          4716 => x"ee",
          4717 => x"51",
          4718 => x"74",
          4719 => x"38",
          4720 => x"08",
          4721 => x"ff",
          4722 => x"74",
          4723 => x"29",
          4724 => x"05",
          4725 => x"82",
          4726 => x"58",
          4727 => x"75",
          4728 => x"fa",
          4729 => x"ee",
          4730 => x"05",
          4731 => x"34",
          4732 => x"08",
          4733 => x"ff",
          4734 => x"82",
          4735 => x"79",
          4736 => x"3f",
          4737 => x"08",
          4738 => x"54",
          4739 => x"82",
          4740 => x"54",
          4741 => x"8f",
          4742 => x"73",
          4743 => x"f1",
          4744 => x"39",
          4745 => x"80",
          4746 => x"9c",
          4747 => x"82",
          4748 => x"79",
          4749 => x"0c",
          4750 => x"04",
          4751 => x"33",
          4752 => x"2e",
          4753 => x"82",
          4754 => x"52",
          4755 => x"9e",
          4756 => x"ee",
          4757 => x"05",
          4758 => x"ee",
          4759 => x"81",
          4760 => x"dd",
          4761 => x"9c",
          4762 => x"98",
          4763 => x"73",
          4764 => x"8c",
          4765 => x"54",
          4766 => x"98",
          4767 => x"2b",
          4768 => x"75",
          4769 => x"56",
          4770 => x"74",
          4771 => x"74",
          4772 => x"14",
          4773 => x"82",
          4774 => x"52",
          4775 => x"ff",
          4776 => x"74",
          4777 => x"29",
          4778 => x"05",
          4779 => x"82",
          4780 => x"58",
          4781 => x"75",
          4782 => x"82",
          4783 => x"52",
          4784 => x"9d",
          4785 => x"ee",
          4786 => x"98",
          4787 => x"2c",
          4788 => x"33",
          4789 => x"57",
          4790 => x"f8",
          4791 => x"f2",
          4792 => x"88",
          4793 => x"cb",
          4794 => x"80",
          4795 => x"80",
          4796 => x"98",
          4797 => x"98",
          4798 => x"55",
          4799 => x"de",
          4800 => x"39",
          4801 => x"33",
          4802 => x"06",
          4803 => x"33",
          4804 => x"74",
          4805 => x"e8",
          4806 => x"bc",
          4807 => x"14",
          4808 => x"ee",
          4809 => x"1a",
          4810 => x"54",
          4811 => x"3f",
          4812 => x"33",
          4813 => x"06",
          4814 => x"33",
          4815 => x"75",
          4816 => x"38",
          4817 => x"82",
          4818 => x"80",
          4819 => x"a0",
          4820 => x"3f",
          4821 => x"ee",
          4822 => x"0b",
          4823 => x"34",
          4824 => x"7a",
          4825 => x"d5",
          4826 => x"74",
          4827 => x"38",
          4828 => x"a5",
          4829 => x"d6",
          4830 => x"ee",
          4831 => x"d6",
          4832 => x"ff",
          4833 => x"53",
          4834 => x"51",
          4835 => x"3f",
          4836 => x"c0",
          4837 => x"29",
          4838 => x"05",
          4839 => x"56",
          4840 => x"2e",
          4841 => x"51",
          4842 => x"3f",
          4843 => x"08",
          4844 => x"34",
          4845 => x"08",
          4846 => x"81",
          4847 => x"52",
          4848 => x"a6",
          4849 => x"1b",
          4850 => x"39",
          4851 => x"74",
          4852 => x"ac",
          4853 => x"ff",
          4854 => x"99",
          4855 => x"2e",
          4856 => x"ae",
          4857 => x"cc",
          4858 => x"80",
          4859 => x"74",
          4860 => x"92",
          4861 => x"d8",
          4862 => x"98",
          4863 => x"d8",
          4864 => x"06",
          4865 => x"74",
          4866 => x"ff",
          4867 => x"80",
          4868 => x"84",
          4869 => x"d0",
          4870 => x"56",
          4871 => x"2e",
          4872 => x"51",
          4873 => x"3f",
          4874 => x"08",
          4875 => x"34",
          4876 => x"08",
          4877 => x"81",
          4878 => x"52",
          4879 => x"a5",
          4880 => x"1b",
          4881 => x"ff",
          4882 => x"39",
          4883 => x"98",
          4884 => x"34",
          4885 => x"53",
          4886 => x"33",
          4887 => x"ec",
          4888 => x"9c",
          4889 => x"9c",
          4890 => x"ff",
          4891 => x"98",
          4892 => x"54",
          4893 => x"f5",
          4894 => x"f2",
          4895 => x"81",
          4896 => x"82",
          4897 => x"74",
          4898 => x"52",
          4899 => x"a3",
          4900 => x"39",
          4901 => x"33",
          4902 => x"2e",
          4903 => x"82",
          4904 => x"52",
          4905 => x"9a",
          4906 => x"ee",
          4907 => x"05",
          4908 => x"ee",
          4909 => x"c8",
          4910 => x"0d",
          4911 => x"33",
          4912 => x"2e",
          4913 => x"a0",
          4914 => x"c4",
          4915 => x"82",
          4916 => x"98",
          4917 => x"c4",
          4918 => x"38",
          4919 => x"d6",
          4920 => x"0b",
          4921 => x"0c",
          4922 => x"08",
          4923 => x"d6",
          4924 => x"70",
          4925 => x"d6",
          4926 => x"87",
          4927 => x"11",
          4928 => x"c0",
          4929 => x"51",
          4930 => x"12",
          4931 => x"82",
          4932 => x"81",
          4933 => x"c8",
          4934 => x"82",
          4935 => x"25",
          4936 => x"d6",
          4937 => x"05",
          4938 => x"0c",
          4939 => x"d6",
          4940 => x"87",
          4941 => x"82",
          4942 => x"80",
          4943 => x"c8",
          4944 => x"82",
          4945 => x"83",
          4946 => x"ff",
          4947 => x"d8",
          4948 => x"3d",
          4949 => x"f4",
          4950 => x"d0",
          4951 => x"0b",
          4952 => x"23",
          4953 => x"80",
          4954 => x"f4",
          4955 => x"a2",
          4956 => x"d0",
          4957 => x"58",
          4958 => x"81",
          4959 => x"15",
          4960 => x"d0",
          4961 => x"84",
          4962 => x"85",
          4963 => x"d6",
          4964 => x"77",
          4965 => x"76",
          4966 => x"82",
          4967 => x"82",
          4968 => x"ff",
          4969 => x"80",
          4970 => x"ff",
          4971 => x"88",
          4972 => x"55",
          4973 => x"17",
          4974 => x"17",
          4975 => x"cc",
          4976 => x"29",
          4977 => x"08",
          4978 => x"51",
          4979 => x"82",
          4980 => x"83",
          4981 => x"3d",
          4982 => x"3d",
          4983 => x"81",
          4984 => x"27",
          4985 => x"12",
          4986 => x"11",
          4987 => x"ff",
          4988 => x"51",
          4989 => x"d8",
          4990 => x"0d",
          4991 => x"0d",
          4992 => x"22",
          4993 => x"aa",
          4994 => x"05",
          4995 => x"08",
          4996 => x"71",
          4997 => x"2b",
          4998 => x"33",
          4999 => x"71",
          5000 => x"02",
          5001 => x"05",
          5002 => x"ff",
          5003 => x"70",
          5004 => x"51",
          5005 => x"5b",
          5006 => x"54",
          5007 => x"34",
          5008 => x"34",
          5009 => x"08",
          5010 => x"2a",
          5011 => x"82",
          5012 => x"83",
          5013 => x"d6",
          5014 => x"17",
          5015 => x"12",
          5016 => x"2b",
          5017 => x"2b",
          5018 => x"06",
          5019 => x"52",
          5020 => x"83",
          5021 => x"70",
          5022 => x"54",
          5023 => x"12",
          5024 => x"ff",
          5025 => x"83",
          5026 => x"d6",
          5027 => x"56",
          5028 => x"72",
          5029 => x"89",
          5030 => x"fb",
          5031 => x"d6",
          5032 => x"84",
          5033 => x"22",
          5034 => x"72",
          5035 => x"33",
          5036 => x"71",
          5037 => x"83",
          5038 => x"5b",
          5039 => x"52",
          5040 => x"12",
          5041 => x"33",
          5042 => x"07",
          5043 => x"54",
          5044 => x"70",
          5045 => x"73",
          5046 => x"82",
          5047 => x"70",
          5048 => x"33",
          5049 => x"71",
          5050 => x"83",
          5051 => x"59",
          5052 => x"05",
          5053 => x"87",
          5054 => x"88",
          5055 => x"88",
          5056 => x"56",
          5057 => x"13",
          5058 => x"13",
          5059 => x"d0",
          5060 => x"33",
          5061 => x"71",
          5062 => x"70",
          5063 => x"06",
          5064 => x"53",
          5065 => x"53",
          5066 => x"70",
          5067 => x"87",
          5068 => x"fa",
          5069 => x"a2",
          5070 => x"d6",
          5071 => x"83",
          5072 => x"70",
          5073 => x"33",
          5074 => x"07",
          5075 => x"15",
          5076 => x"12",
          5077 => x"2b",
          5078 => x"07",
          5079 => x"55",
          5080 => x"57",
          5081 => x"80",
          5082 => x"38",
          5083 => x"ab",
          5084 => x"d0",
          5085 => x"70",
          5086 => x"33",
          5087 => x"71",
          5088 => x"74",
          5089 => x"81",
          5090 => x"88",
          5091 => x"83",
          5092 => x"f8",
          5093 => x"54",
          5094 => x"58",
          5095 => x"74",
          5096 => x"52",
          5097 => x"34",
          5098 => x"34",
          5099 => x"08",
          5100 => x"33",
          5101 => x"71",
          5102 => x"83",
          5103 => x"59",
          5104 => x"05",
          5105 => x"12",
          5106 => x"2b",
          5107 => x"ff",
          5108 => x"88",
          5109 => x"52",
          5110 => x"74",
          5111 => x"15",
          5112 => x"0d",
          5113 => x"0d",
          5114 => x"08",
          5115 => x"9e",
          5116 => x"83",
          5117 => x"82",
          5118 => x"12",
          5119 => x"2b",
          5120 => x"07",
          5121 => x"52",
          5122 => x"05",
          5123 => x"13",
          5124 => x"2b",
          5125 => x"05",
          5126 => x"71",
          5127 => x"2a",
          5128 => x"53",
          5129 => x"34",
          5130 => x"34",
          5131 => x"08",
          5132 => x"33",
          5133 => x"71",
          5134 => x"83",
          5135 => x"59",
          5136 => x"05",
          5137 => x"83",
          5138 => x"88",
          5139 => x"88",
          5140 => x"56",
          5141 => x"13",
          5142 => x"13",
          5143 => x"d0",
          5144 => x"11",
          5145 => x"33",
          5146 => x"07",
          5147 => x"0c",
          5148 => x"3d",
          5149 => x"3d",
          5150 => x"d6",
          5151 => x"83",
          5152 => x"ff",
          5153 => x"53",
          5154 => x"a7",
          5155 => x"d0",
          5156 => x"2b",
          5157 => x"11",
          5158 => x"33",
          5159 => x"71",
          5160 => x"75",
          5161 => x"81",
          5162 => x"98",
          5163 => x"2b",
          5164 => x"40",
          5165 => x"58",
          5166 => x"72",
          5167 => x"38",
          5168 => x"52",
          5169 => x"9d",
          5170 => x"39",
          5171 => x"85",
          5172 => x"8b",
          5173 => x"2b",
          5174 => x"79",
          5175 => x"51",
          5176 => x"76",
          5177 => x"75",
          5178 => x"56",
          5179 => x"34",
          5180 => x"08",
          5181 => x"12",
          5182 => x"33",
          5183 => x"07",
          5184 => x"54",
          5185 => x"53",
          5186 => x"34",
          5187 => x"34",
          5188 => x"08",
          5189 => x"0b",
          5190 => x"80",
          5191 => x"34",
          5192 => x"08",
          5193 => x"14",
          5194 => x"14",
          5195 => x"d0",
          5196 => x"33",
          5197 => x"71",
          5198 => x"70",
          5199 => x"07",
          5200 => x"53",
          5201 => x"54",
          5202 => x"72",
          5203 => x"8b",
          5204 => x"ff",
          5205 => x"52",
          5206 => x"08",
          5207 => x"f2",
          5208 => x"2e",
          5209 => x"51",
          5210 => x"83",
          5211 => x"f5",
          5212 => x"7e",
          5213 => x"e2",
          5214 => x"d8",
          5215 => x"ff",
          5216 => x"d0",
          5217 => x"33",
          5218 => x"71",
          5219 => x"70",
          5220 => x"58",
          5221 => x"ff",
          5222 => x"2e",
          5223 => x"75",
          5224 => x"70",
          5225 => x"33",
          5226 => x"07",
          5227 => x"ff",
          5228 => x"70",
          5229 => x"06",
          5230 => x"52",
          5231 => x"59",
          5232 => x"27",
          5233 => x"80",
          5234 => x"75",
          5235 => x"84",
          5236 => x"16",
          5237 => x"2b",
          5238 => x"75",
          5239 => x"81",
          5240 => x"85",
          5241 => x"59",
          5242 => x"83",
          5243 => x"d0",
          5244 => x"33",
          5245 => x"71",
          5246 => x"70",
          5247 => x"06",
          5248 => x"56",
          5249 => x"75",
          5250 => x"81",
          5251 => x"79",
          5252 => x"cc",
          5253 => x"74",
          5254 => x"c4",
          5255 => x"2e",
          5256 => x"89",
          5257 => x"f8",
          5258 => x"ac",
          5259 => x"80",
          5260 => x"75",
          5261 => x"3f",
          5262 => x"08",
          5263 => x"11",
          5264 => x"33",
          5265 => x"71",
          5266 => x"53",
          5267 => x"74",
          5268 => x"70",
          5269 => x"06",
          5270 => x"5c",
          5271 => x"78",
          5272 => x"76",
          5273 => x"57",
          5274 => x"34",
          5275 => x"08",
          5276 => x"71",
          5277 => x"86",
          5278 => x"12",
          5279 => x"2b",
          5280 => x"2a",
          5281 => x"53",
          5282 => x"73",
          5283 => x"75",
          5284 => x"82",
          5285 => x"70",
          5286 => x"33",
          5287 => x"71",
          5288 => x"83",
          5289 => x"5d",
          5290 => x"05",
          5291 => x"15",
          5292 => x"15",
          5293 => x"d0",
          5294 => x"71",
          5295 => x"33",
          5296 => x"71",
          5297 => x"70",
          5298 => x"5a",
          5299 => x"54",
          5300 => x"34",
          5301 => x"34",
          5302 => x"08",
          5303 => x"54",
          5304 => x"d8",
          5305 => x"0d",
          5306 => x"0d",
          5307 => x"d6",
          5308 => x"38",
          5309 => x"71",
          5310 => x"2e",
          5311 => x"51",
          5312 => x"82",
          5313 => x"53",
          5314 => x"d8",
          5315 => x"0d",
          5316 => x"0d",
          5317 => x"5c",
          5318 => x"40",
          5319 => x"08",
          5320 => x"81",
          5321 => x"f4",
          5322 => x"8e",
          5323 => x"ff",
          5324 => x"d6",
          5325 => x"83",
          5326 => x"8b",
          5327 => x"fc",
          5328 => x"54",
          5329 => x"7e",
          5330 => x"3f",
          5331 => x"08",
          5332 => x"06",
          5333 => x"08",
          5334 => x"83",
          5335 => x"ff",
          5336 => x"83",
          5337 => x"70",
          5338 => x"33",
          5339 => x"07",
          5340 => x"70",
          5341 => x"06",
          5342 => x"fc",
          5343 => x"29",
          5344 => x"81",
          5345 => x"88",
          5346 => x"90",
          5347 => x"4e",
          5348 => x"52",
          5349 => x"41",
          5350 => x"5b",
          5351 => x"8f",
          5352 => x"ff",
          5353 => x"31",
          5354 => x"ff",
          5355 => x"82",
          5356 => x"17",
          5357 => x"2b",
          5358 => x"29",
          5359 => x"81",
          5360 => x"98",
          5361 => x"2b",
          5362 => x"45",
          5363 => x"73",
          5364 => x"38",
          5365 => x"70",
          5366 => x"06",
          5367 => x"7b",
          5368 => x"38",
          5369 => x"73",
          5370 => x"81",
          5371 => x"78",
          5372 => x"3f",
          5373 => x"ff",
          5374 => x"e5",
          5375 => x"38",
          5376 => x"89",
          5377 => x"f6",
          5378 => x"a5",
          5379 => x"55",
          5380 => x"80",
          5381 => x"1d",
          5382 => x"83",
          5383 => x"88",
          5384 => x"57",
          5385 => x"3f",
          5386 => x"51",
          5387 => x"82",
          5388 => x"83",
          5389 => x"7e",
          5390 => x"70",
          5391 => x"d6",
          5392 => x"84",
          5393 => x"59",
          5394 => x"3f",
          5395 => x"08",
          5396 => x"75",
          5397 => x"06",
          5398 => x"85",
          5399 => x"54",
          5400 => x"80",
          5401 => x"51",
          5402 => x"82",
          5403 => x"1d",
          5404 => x"83",
          5405 => x"88",
          5406 => x"43",
          5407 => x"3f",
          5408 => x"51",
          5409 => x"82",
          5410 => x"83",
          5411 => x"7e",
          5412 => x"70",
          5413 => x"d6",
          5414 => x"84",
          5415 => x"59",
          5416 => x"3f",
          5417 => x"08",
          5418 => x"60",
          5419 => x"55",
          5420 => x"ff",
          5421 => x"a9",
          5422 => x"52",
          5423 => x"3f",
          5424 => x"08",
          5425 => x"d8",
          5426 => x"93",
          5427 => x"73",
          5428 => x"d8",
          5429 => x"94",
          5430 => x"51",
          5431 => x"7a",
          5432 => x"27",
          5433 => x"53",
          5434 => x"51",
          5435 => x"7a",
          5436 => x"82",
          5437 => x"05",
          5438 => x"f6",
          5439 => x"54",
          5440 => x"d8",
          5441 => x"0d",
          5442 => x"0d",
          5443 => x"70",
          5444 => x"d5",
          5445 => x"d8",
          5446 => x"d6",
          5447 => x"2e",
          5448 => x"53",
          5449 => x"d6",
          5450 => x"ff",
          5451 => x"74",
          5452 => x"0c",
          5453 => x"04",
          5454 => x"02",
          5455 => x"51",
          5456 => x"72",
          5457 => x"82",
          5458 => x"33",
          5459 => x"d6",
          5460 => x"3d",
          5461 => x"3d",
          5462 => x"05",
          5463 => x"05",
          5464 => x"56",
          5465 => x"72",
          5466 => x"e0",
          5467 => x"2b",
          5468 => x"8c",
          5469 => x"88",
          5470 => x"2e",
          5471 => x"88",
          5472 => x"0c",
          5473 => x"8c",
          5474 => x"71",
          5475 => x"87",
          5476 => x"0c",
          5477 => x"08",
          5478 => x"51",
          5479 => x"2e",
          5480 => x"c0",
          5481 => x"51",
          5482 => x"71",
          5483 => x"80",
          5484 => x"92",
          5485 => x"98",
          5486 => x"70",
          5487 => x"38",
          5488 => x"d4",
          5489 => x"d6",
          5490 => x"51",
          5491 => x"d8",
          5492 => x"0d",
          5493 => x"0d",
          5494 => x"02",
          5495 => x"05",
          5496 => x"58",
          5497 => x"52",
          5498 => x"3f",
          5499 => x"08",
          5500 => x"54",
          5501 => x"be",
          5502 => x"75",
          5503 => x"c0",
          5504 => x"87",
          5505 => x"12",
          5506 => x"84",
          5507 => x"40",
          5508 => x"85",
          5509 => x"98",
          5510 => x"7d",
          5511 => x"0c",
          5512 => x"85",
          5513 => x"06",
          5514 => x"71",
          5515 => x"38",
          5516 => x"71",
          5517 => x"05",
          5518 => x"19",
          5519 => x"a2",
          5520 => x"71",
          5521 => x"38",
          5522 => x"83",
          5523 => x"38",
          5524 => x"8a",
          5525 => x"98",
          5526 => x"71",
          5527 => x"c0",
          5528 => x"52",
          5529 => x"87",
          5530 => x"80",
          5531 => x"81",
          5532 => x"c0",
          5533 => x"53",
          5534 => x"82",
          5535 => x"71",
          5536 => x"1a",
          5537 => x"84",
          5538 => x"19",
          5539 => x"06",
          5540 => x"79",
          5541 => x"38",
          5542 => x"80",
          5543 => x"87",
          5544 => x"26",
          5545 => x"73",
          5546 => x"06",
          5547 => x"2e",
          5548 => x"52",
          5549 => x"82",
          5550 => x"8f",
          5551 => x"f3",
          5552 => x"62",
          5553 => x"05",
          5554 => x"57",
          5555 => x"83",
          5556 => x"52",
          5557 => x"3f",
          5558 => x"08",
          5559 => x"54",
          5560 => x"2e",
          5561 => x"81",
          5562 => x"74",
          5563 => x"c0",
          5564 => x"87",
          5565 => x"12",
          5566 => x"84",
          5567 => x"5f",
          5568 => x"0b",
          5569 => x"8c",
          5570 => x"0c",
          5571 => x"80",
          5572 => x"70",
          5573 => x"81",
          5574 => x"54",
          5575 => x"8c",
          5576 => x"81",
          5577 => x"7c",
          5578 => x"58",
          5579 => x"70",
          5580 => x"52",
          5581 => x"8a",
          5582 => x"98",
          5583 => x"71",
          5584 => x"c0",
          5585 => x"52",
          5586 => x"87",
          5587 => x"80",
          5588 => x"81",
          5589 => x"c0",
          5590 => x"53",
          5591 => x"82",
          5592 => x"71",
          5593 => x"19",
          5594 => x"81",
          5595 => x"ff",
          5596 => x"19",
          5597 => x"78",
          5598 => x"38",
          5599 => x"80",
          5600 => x"87",
          5601 => x"26",
          5602 => x"73",
          5603 => x"06",
          5604 => x"2e",
          5605 => x"52",
          5606 => x"82",
          5607 => x"8f",
          5608 => x"fa",
          5609 => x"02",
          5610 => x"05",
          5611 => x"05",
          5612 => x"71",
          5613 => x"57",
          5614 => x"82",
          5615 => x"81",
          5616 => x"54",
          5617 => x"38",
          5618 => x"c0",
          5619 => x"81",
          5620 => x"2e",
          5621 => x"71",
          5622 => x"38",
          5623 => x"87",
          5624 => x"11",
          5625 => x"80",
          5626 => x"80",
          5627 => x"83",
          5628 => x"38",
          5629 => x"72",
          5630 => x"2a",
          5631 => x"51",
          5632 => x"80",
          5633 => x"87",
          5634 => x"08",
          5635 => x"38",
          5636 => x"8c",
          5637 => x"96",
          5638 => x"0c",
          5639 => x"8c",
          5640 => x"08",
          5641 => x"51",
          5642 => x"38",
          5643 => x"56",
          5644 => x"80",
          5645 => x"85",
          5646 => x"77",
          5647 => x"83",
          5648 => x"75",
          5649 => x"d6",
          5650 => x"3d",
          5651 => x"3d",
          5652 => x"11",
          5653 => x"71",
          5654 => x"82",
          5655 => x"53",
          5656 => x"0d",
          5657 => x"0d",
          5658 => x"33",
          5659 => x"71",
          5660 => x"88",
          5661 => x"14",
          5662 => x"07",
          5663 => x"33",
          5664 => x"d6",
          5665 => x"53",
          5666 => x"52",
          5667 => x"04",
          5668 => x"73",
          5669 => x"92",
          5670 => x"52",
          5671 => x"81",
          5672 => x"70",
          5673 => x"70",
          5674 => x"3d",
          5675 => x"3d",
          5676 => x"52",
          5677 => x"70",
          5678 => x"34",
          5679 => x"51",
          5680 => x"81",
          5681 => x"70",
          5682 => x"70",
          5683 => x"05",
          5684 => x"88",
          5685 => x"72",
          5686 => x"0d",
          5687 => x"0d",
          5688 => x"54",
          5689 => x"80",
          5690 => x"71",
          5691 => x"53",
          5692 => x"81",
          5693 => x"ff",
          5694 => x"39",
          5695 => x"04",
          5696 => x"75",
          5697 => x"52",
          5698 => x"70",
          5699 => x"34",
          5700 => x"70",
          5701 => x"3d",
          5702 => x"3d",
          5703 => x"79",
          5704 => x"74",
          5705 => x"56",
          5706 => x"81",
          5707 => x"71",
          5708 => x"16",
          5709 => x"52",
          5710 => x"86",
          5711 => x"2e",
          5712 => x"82",
          5713 => x"86",
          5714 => x"fe",
          5715 => x"76",
          5716 => x"39",
          5717 => x"8a",
          5718 => x"51",
          5719 => x"71",
          5720 => x"33",
          5721 => x"0c",
          5722 => x"04",
          5723 => x"d6",
          5724 => x"fb",
          5725 => x"70",
          5726 => x"81",
          5727 => x"70",
          5728 => x"56",
          5729 => x"55",
          5730 => x"08",
          5731 => x"80",
          5732 => x"83",
          5733 => x"51",
          5734 => x"3f",
          5735 => x"08",
          5736 => x"06",
          5737 => x"2e",
          5738 => x"76",
          5739 => x"74",
          5740 => x"0c",
          5741 => x"04",
          5742 => x"7b",
          5743 => x"83",
          5744 => x"5a",
          5745 => x"80",
          5746 => x"54",
          5747 => x"53",
          5748 => x"53",
          5749 => x"52",
          5750 => x"3f",
          5751 => x"08",
          5752 => x"81",
          5753 => x"82",
          5754 => x"83",
          5755 => x"16",
          5756 => x"18",
          5757 => x"18",
          5758 => x"58",
          5759 => x"9f",
          5760 => x"33",
          5761 => x"2e",
          5762 => x"93",
          5763 => x"76",
          5764 => x"52",
          5765 => x"51",
          5766 => x"83",
          5767 => x"79",
          5768 => x"0c",
          5769 => x"04",
          5770 => x"78",
          5771 => x"80",
          5772 => x"17",
          5773 => x"38",
          5774 => x"fc",
          5775 => x"d8",
          5776 => x"d6",
          5777 => x"38",
          5778 => x"53",
          5779 => x"81",
          5780 => x"f7",
          5781 => x"d6",
          5782 => x"2e",
          5783 => x"55",
          5784 => x"b4",
          5785 => x"82",
          5786 => x"88",
          5787 => x"f8",
          5788 => x"70",
          5789 => x"c0",
          5790 => x"d8",
          5791 => x"d6",
          5792 => x"91",
          5793 => x"55",
          5794 => x"09",
          5795 => x"f0",
          5796 => x"33",
          5797 => x"2e",
          5798 => x"80",
          5799 => x"80",
          5800 => x"d8",
          5801 => x"17",
          5802 => x"fc",
          5803 => x"d4",
          5804 => x"b6",
          5805 => x"d8",
          5806 => x"85",
          5807 => x"75",
          5808 => x"3f",
          5809 => x"e4",
          5810 => x"9c",
          5811 => x"de",
          5812 => x"08",
          5813 => x"17",
          5814 => x"3f",
          5815 => x"52",
          5816 => x"51",
          5817 => x"a4",
          5818 => x"05",
          5819 => x"0c",
          5820 => x"75",
          5821 => x"33",
          5822 => x"3f",
          5823 => x"34",
          5824 => x"52",
          5825 => x"51",
          5826 => x"82",
          5827 => x"80",
          5828 => x"81",
          5829 => x"d6",
          5830 => x"3d",
          5831 => x"3d",
          5832 => x"1a",
          5833 => x"fe",
          5834 => x"54",
          5835 => x"73",
          5836 => x"8a",
          5837 => x"71",
          5838 => x"08",
          5839 => x"75",
          5840 => x"0c",
          5841 => x"04",
          5842 => x"7a",
          5843 => x"56",
          5844 => x"77",
          5845 => x"38",
          5846 => x"08",
          5847 => x"38",
          5848 => x"54",
          5849 => x"2e",
          5850 => x"72",
          5851 => x"38",
          5852 => x"8d",
          5853 => x"39",
          5854 => x"81",
          5855 => x"b6",
          5856 => x"2a",
          5857 => x"2a",
          5858 => x"05",
          5859 => x"55",
          5860 => x"82",
          5861 => x"81",
          5862 => x"83",
          5863 => x"b8",
          5864 => x"17",
          5865 => x"a8",
          5866 => x"55",
          5867 => x"57",
          5868 => x"3f",
          5869 => x"08",
          5870 => x"74",
          5871 => x"14",
          5872 => x"70",
          5873 => x"07",
          5874 => x"71",
          5875 => x"52",
          5876 => x"72",
          5877 => x"75",
          5878 => x"58",
          5879 => x"76",
          5880 => x"15",
          5881 => x"73",
          5882 => x"3f",
          5883 => x"08",
          5884 => x"76",
          5885 => x"06",
          5886 => x"05",
          5887 => x"3f",
          5888 => x"08",
          5889 => x"06",
          5890 => x"76",
          5891 => x"15",
          5892 => x"73",
          5893 => x"3f",
          5894 => x"08",
          5895 => x"82",
          5896 => x"06",
          5897 => x"05",
          5898 => x"3f",
          5899 => x"08",
          5900 => x"58",
          5901 => x"58",
          5902 => x"d8",
          5903 => x"0d",
          5904 => x"0d",
          5905 => x"5a",
          5906 => x"59",
          5907 => x"82",
          5908 => x"9c",
          5909 => x"82",
          5910 => x"33",
          5911 => x"2e",
          5912 => x"72",
          5913 => x"38",
          5914 => x"8d",
          5915 => x"39",
          5916 => x"81",
          5917 => x"f7",
          5918 => x"2a",
          5919 => x"2a",
          5920 => x"05",
          5921 => x"55",
          5922 => x"82",
          5923 => x"59",
          5924 => x"08",
          5925 => x"74",
          5926 => x"16",
          5927 => x"16",
          5928 => x"59",
          5929 => x"53",
          5930 => x"8f",
          5931 => x"2b",
          5932 => x"74",
          5933 => x"71",
          5934 => x"72",
          5935 => x"0b",
          5936 => x"74",
          5937 => x"17",
          5938 => x"75",
          5939 => x"3f",
          5940 => x"08",
          5941 => x"d8",
          5942 => x"38",
          5943 => x"06",
          5944 => x"78",
          5945 => x"54",
          5946 => x"77",
          5947 => x"33",
          5948 => x"71",
          5949 => x"51",
          5950 => x"34",
          5951 => x"76",
          5952 => x"17",
          5953 => x"75",
          5954 => x"3f",
          5955 => x"08",
          5956 => x"d8",
          5957 => x"38",
          5958 => x"ff",
          5959 => x"10",
          5960 => x"76",
          5961 => x"51",
          5962 => x"be",
          5963 => x"2a",
          5964 => x"05",
          5965 => x"f9",
          5966 => x"d6",
          5967 => x"82",
          5968 => x"ab",
          5969 => x"0a",
          5970 => x"2b",
          5971 => x"70",
          5972 => x"70",
          5973 => x"54",
          5974 => x"82",
          5975 => x"8f",
          5976 => x"07",
          5977 => x"f6",
          5978 => x"0b",
          5979 => x"78",
          5980 => x"0c",
          5981 => x"04",
          5982 => x"7a",
          5983 => x"08",
          5984 => x"59",
          5985 => x"a4",
          5986 => x"17",
          5987 => x"38",
          5988 => x"aa",
          5989 => x"73",
          5990 => x"fd",
          5991 => x"d6",
          5992 => x"82",
          5993 => x"80",
          5994 => x"39",
          5995 => x"eb",
          5996 => x"80",
          5997 => x"d6",
          5998 => x"80",
          5999 => x"52",
          6000 => x"84",
          6001 => x"d8",
          6002 => x"d6",
          6003 => x"2e",
          6004 => x"82",
          6005 => x"81",
          6006 => x"82",
          6007 => x"ff",
          6008 => x"80",
          6009 => x"75",
          6010 => x"3f",
          6011 => x"08",
          6012 => x"16",
          6013 => x"94",
          6014 => x"55",
          6015 => x"27",
          6016 => x"15",
          6017 => x"84",
          6018 => x"07",
          6019 => x"17",
          6020 => x"76",
          6021 => x"a6",
          6022 => x"73",
          6023 => x"0c",
          6024 => x"04",
          6025 => x"7c",
          6026 => x"59",
          6027 => x"95",
          6028 => x"08",
          6029 => x"2e",
          6030 => x"17",
          6031 => x"b2",
          6032 => x"ae",
          6033 => x"7a",
          6034 => x"3f",
          6035 => x"82",
          6036 => x"27",
          6037 => x"82",
          6038 => x"55",
          6039 => x"08",
          6040 => x"d2",
          6041 => x"08",
          6042 => x"08",
          6043 => x"38",
          6044 => x"17",
          6045 => x"54",
          6046 => x"82",
          6047 => x"7a",
          6048 => x"06",
          6049 => x"81",
          6050 => x"17",
          6051 => x"83",
          6052 => x"75",
          6053 => x"f9",
          6054 => x"59",
          6055 => x"08",
          6056 => x"81",
          6057 => x"82",
          6058 => x"59",
          6059 => x"08",
          6060 => x"70",
          6061 => x"25",
          6062 => x"82",
          6063 => x"54",
          6064 => x"55",
          6065 => x"38",
          6066 => x"08",
          6067 => x"38",
          6068 => x"54",
          6069 => x"90",
          6070 => x"18",
          6071 => x"38",
          6072 => x"39",
          6073 => x"38",
          6074 => x"16",
          6075 => x"08",
          6076 => x"38",
          6077 => x"78",
          6078 => x"38",
          6079 => x"51",
          6080 => x"82",
          6081 => x"80",
          6082 => x"80",
          6083 => x"d8",
          6084 => x"09",
          6085 => x"38",
          6086 => x"08",
          6087 => x"d8",
          6088 => x"30",
          6089 => x"80",
          6090 => x"07",
          6091 => x"55",
          6092 => x"38",
          6093 => x"09",
          6094 => x"ae",
          6095 => x"80",
          6096 => x"53",
          6097 => x"51",
          6098 => x"82",
          6099 => x"82",
          6100 => x"30",
          6101 => x"d8",
          6102 => x"25",
          6103 => x"79",
          6104 => x"38",
          6105 => x"8f",
          6106 => x"79",
          6107 => x"f9",
          6108 => x"d6",
          6109 => x"74",
          6110 => x"90",
          6111 => x"17",
          6112 => x"94",
          6113 => x"54",
          6114 => x"86",
          6115 => x"94",
          6116 => x"17",
          6117 => x"54",
          6118 => x"34",
          6119 => x"56",
          6120 => x"90",
          6121 => x"80",
          6122 => x"82",
          6123 => x"55",
          6124 => x"56",
          6125 => x"82",
          6126 => x"8c",
          6127 => x"f8",
          6128 => x"70",
          6129 => x"f0",
          6130 => x"d8",
          6131 => x"56",
          6132 => x"08",
          6133 => x"7b",
          6134 => x"f6",
          6135 => x"d6",
          6136 => x"d6",
          6137 => x"17",
          6138 => x"80",
          6139 => x"b8",
          6140 => x"57",
          6141 => x"77",
          6142 => x"81",
          6143 => x"15",
          6144 => x"78",
          6145 => x"81",
          6146 => x"53",
          6147 => x"15",
          6148 => x"ab",
          6149 => x"d8",
          6150 => x"df",
          6151 => x"22",
          6152 => x"30",
          6153 => x"70",
          6154 => x"51",
          6155 => x"82",
          6156 => x"8a",
          6157 => x"f8",
          6158 => x"7c",
          6159 => x"56",
          6160 => x"80",
          6161 => x"f1",
          6162 => x"06",
          6163 => x"e9",
          6164 => x"18",
          6165 => x"08",
          6166 => x"38",
          6167 => x"82",
          6168 => x"38",
          6169 => x"54",
          6170 => x"74",
          6171 => x"82",
          6172 => x"22",
          6173 => x"79",
          6174 => x"38",
          6175 => x"98",
          6176 => x"cd",
          6177 => x"22",
          6178 => x"54",
          6179 => x"26",
          6180 => x"52",
          6181 => x"b0",
          6182 => x"d8",
          6183 => x"d6",
          6184 => x"2e",
          6185 => x"0b",
          6186 => x"08",
          6187 => x"9c",
          6188 => x"d6",
          6189 => x"85",
          6190 => x"bd",
          6191 => x"31",
          6192 => x"73",
          6193 => x"f4",
          6194 => x"d6",
          6195 => x"18",
          6196 => x"18",
          6197 => x"08",
          6198 => x"72",
          6199 => x"38",
          6200 => x"58",
          6201 => x"89",
          6202 => x"18",
          6203 => x"ff",
          6204 => x"05",
          6205 => x"80",
          6206 => x"d6",
          6207 => x"3d",
          6208 => x"3d",
          6209 => x"08",
          6210 => x"a0",
          6211 => x"54",
          6212 => x"77",
          6213 => x"80",
          6214 => x"0c",
          6215 => x"53",
          6216 => x"80",
          6217 => x"38",
          6218 => x"06",
          6219 => x"b5",
          6220 => x"98",
          6221 => x"14",
          6222 => x"92",
          6223 => x"2a",
          6224 => x"56",
          6225 => x"26",
          6226 => x"80",
          6227 => x"16",
          6228 => x"77",
          6229 => x"53",
          6230 => x"38",
          6231 => x"51",
          6232 => x"82",
          6233 => x"53",
          6234 => x"0b",
          6235 => x"08",
          6236 => x"38",
          6237 => x"d6",
          6238 => x"2e",
          6239 => x"9c",
          6240 => x"d6",
          6241 => x"80",
          6242 => x"8a",
          6243 => x"15",
          6244 => x"80",
          6245 => x"14",
          6246 => x"51",
          6247 => x"82",
          6248 => x"53",
          6249 => x"d6",
          6250 => x"2e",
          6251 => x"82",
          6252 => x"d8",
          6253 => x"ba",
          6254 => x"82",
          6255 => x"ff",
          6256 => x"82",
          6257 => x"52",
          6258 => x"f3",
          6259 => x"d8",
          6260 => x"72",
          6261 => x"72",
          6262 => x"f2",
          6263 => x"d6",
          6264 => x"15",
          6265 => x"15",
          6266 => x"b8",
          6267 => x"0c",
          6268 => x"82",
          6269 => x"8a",
          6270 => x"f7",
          6271 => x"7d",
          6272 => x"5b",
          6273 => x"76",
          6274 => x"3f",
          6275 => x"08",
          6276 => x"d8",
          6277 => x"38",
          6278 => x"08",
          6279 => x"08",
          6280 => x"f0",
          6281 => x"d6",
          6282 => x"82",
          6283 => x"80",
          6284 => x"d6",
          6285 => x"18",
          6286 => x"51",
          6287 => x"81",
          6288 => x"81",
          6289 => x"81",
          6290 => x"d8",
          6291 => x"83",
          6292 => x"77",
          6293 => x"72",
          6294 => x"38",
          6295 => x"75",
          6296 => x"81",
          6297 => x"a5",
          6298 => x"d8",
          6299 => x"52",
          6300 => x"8e",
          6301 => x"d8",
          6302 => x"d6",
          6303 => x"2e",
          6304 => x"73",
          6305 => x"81",
          6306 => x"87",
          6307 => x"d6",
          6308 => x"3d",
          6309 => x"3d",
          6310 => x"11",
          6311 => x"ae",
          6312 => x"d8",
          6313 => x"ff",
          6314 => x"33",
          6315 => x"71",
          6316 => x"81",
          6317 => x"94",
          6318 => x"92",
          6319 => x"d8",
          6320 => x"73",
          6321 => x"82",
          6322 => x"85",
          6323 => x"fc",
          6324 => x"79",
          6325 => x"ff",
          6326 => x"12",
          6327 => x"eb",
          6328 => x"70",
          6329 => x"72",
          6330 => x"81",
          6331 => x"73",
          6332 => x"94",
          6333 => x"98",
          6334 => x"0d",
          6335 => x"0d",
          6336 => x"51",
          6337 => x"81",
          6338 => x"80",
          6339 => x"70",
          6340 => x"33",
          6341 => x"81",
          6342 => x"16",
          6343 => x"51",
          6344 => x"70",
          6345 => x"0c",
          6346 => x"04",
          6347 => x"60",
          6348 => x"84",
          6349 => x"5b",
          6350 => x"5d",
          6351 => x"08",
          6352 => x"80",
          6353 => x"08",
          6354 => x"ed",
          6355 => x"d6",
          6356 => x"82",
          6357 => x"82",
          6358 => x"19",
          6359 => x"55",
          6360 => x"38",
          6361 => x"dc",
          6362 => x"33",
          6363 => x"81",
          6364 => x"53",
          6365 => x"34",
          6366 => x"08",
          6367 => x"e5",
          6368 => x"06",
          6369 => x"56",
          6370 => x"08",
          6371 => x"2e",
          6372 => x"83",
          6373 => x"75",
          6374 => x"72",
          6375 => x"d6",
          6376 => x"df",
          6377 => x"72",
          6378 => x"81",
          6379 => x"81",
          6380 => x"2e",
          6381 => x"ff",
          6382 => x"39",
          6383 => x"09",
          6384 => x"ca",
          6385 => x"2a",
          6386 => x"51",
          6387 => x"2e",
          6388 => x"15",
          6389 => x"bf",
          6390 => x"1c",
          6391 => x"0c",
          6392 => x"73",
          6393 => x"81",
          6394 => x"38",
          6395 => x"53",
          6396 => x"09",
          6397 => x"8f",
          6398 => x"08",
          6399 => x"5a",
          6400 => x"82",
          6401 => x"83",
          6402 => x"53",
          6403 => x"38",
          6404 => x"81",
          6405 => x"29",
          6406 => x"54",
          6407 => x"58",
          6408 => x"17",
          6409 => x"51",
          6410 => x"82",
          6411 => x"83",
          6412 => x"56",
          6413 => x"96",
          6414 => x"fe",
          6415 => x"38",
          6416 => x"76",
          6417 => x"73",
          6418 => x"54",
          6419 => x"83",
          6420 => x"09",
          6421 => x"38",
          6422 => x"8c",
          6423 => x"38",
          6424 => x"86",
          6425 => x"06",
          6426 => x"72",
          6427 => x"38",
          6428 => x"26",
          6429 => x"10",
          6430 => x"73",
          6431 => x"70",
          6432 => x"51",
          6433 => x"81",
          6434 => x"5c",
          6435 => x"93",
          6436 => x"fc",
          6437 => x"d6",
          6438 => x"ff",
          6439 => x"7d",
          6440 => x"ff",
          6441 => x"0c",
          6442 => x"52",
          6443 => x"d2",
          6444 => x"d8",
          6445 => x"d6",
          6446 => x"38",
          6447 => x"fd",
          6448 => x"39",
          6449 => x"1a",
          6450 => x"d6",
          6451 => x"3d",
          6452 => x"3d",
          6453 => x"08",
          6454 => x"52",
          6455 => x"d7",
          6456 => x"d8",
          6457 => x"d6",
          6458 => x"a4",
          6459 => x"70",
          6460 => x"0b",
          6461 => x"98",
          6462 => x"7e",
          6463 => x"3f",
          6464 => x"08",
          6465 => x"d8",
          6466 => x"38",
          6467 => x"70",
          6468 => x"75",
          6469 => x"58",
          6470 => x"8b",
          6471 => x"06",
          6472 => x"06",
          6473 => x"86",
          6474 => x"81",
          6475 => x"c3",
          6476 => x"2a",
          6477 => x"51",
          6478 => x"2e",
          6479 => x"82",
          6480 => x"8f",
          6481 => x"06",
          6482 => x"ab",
          6483 => x"86",
          6484 => x"06",
          6485 => x"73",
          6486 => x"75",
          6487 => x"81",
          6488 => x"73",
          6489 => x"38",
          6490 => x"76",
          6491 => x"70",
          6492 => x"ac",
          6493 => x"5d",
          6494 => x"2e",
          6495 => x"81",
          6496 => x"17",
          6497 => x"76",
          6498 => x"06",
          6499 => x"8c",
          6500 => x"18",
          6501 => x"b6",
          6502 => x"d8",
          6503 => x"ff",
          6504 => x"81",
          6505 => x"33",
          6506 => x"8d",
          6507 => x"59",
          6508 => x"5c",
          6509 => x"d4",
          6510 => x"05",
          6511 => x"3f",
          6512 => x"08",
          6513 => x"06",
          6514 => x"2e",
          6515 => x"81",
          6516 => x"e6",
          6517 => x"80",
          6518 => x"82",
          6519 => x"78",
          6520 => x"22",
          6521 => x"19",
          6522 => x"df",
          6523 => x"82",
          6524 => x"2e",
          6525 => x"80",
          6526 => x"5a",
          6527 => x"83",
          6528 => x"09",
          6529 => x"38",
          6530 => x"8c",
          6531 => x"a5",
          6532 => x"70",
          6533 => x"81",
          6534 => x"57",
          6535 => x"90",
          6536 => x"2e",
          6537 => x"10",
          6538 => x"51",
          6539 => x"38",
          6540 => x"81",
          6541 => x"54",
          6542 => x"ff",
          6543 => x"bb",
          6544 => x"38",
          6545 => x"b5",
          6546 => x"d8",
          6547 => x"06",
          6548 => x"2e",
          6549 => x"19",
          6550 => x"54",
          6551 => x"8b",
          6552 => x"52",
          6553 => x"51",
          6554 => x"82",
          6555 => x"80",
          6556 => x"81",
          6557 => x"0b",
          6558 => x"80",
          6559 => x"f5",
          6560 => x"d6",
          6561 => x"82",
          6562 => x"80",
          6563 => x"38",
          6564 => x"d8",
          6565 => x"0d",
          6566 => x"0d",
          6567 => x"ab",
          6568 => x"a0",
          6569 => x"5a",
          6570 => x"85",
          6571 => x"8c",
          6572 => x"22",
          6573 => x"73",
          6574 => x"38",
          6575 => x"10",
          6576 => x"51",
          6577 => x"39",
          6578 => x"1a",
          6579 => x"3d",
          6580 => x"59",
          6581 => x"02",
          6582 => x"33",
          6583 => x"73",
          6584 => x"a8",
          6585 => x"0b",
          6586 => x"81",
          6587 => x"08",
          6588 => x"8b",
          6589 => x"78",
          6590 => x"3f",
          6591 => x"80",
          6592 => x"56",
          6593 => x"83",
          6594 => x"55",
          6595 => x"2e",
          6596 => x"83",
          6597 => x"82",
          6598 => x"8f",
          6599 => x"06",
          6600 => x"75",
          6601 => x"90",
          6602 => x"06",
          6603 => x"56",
          6604 => x"87",
          6605 => x"a0",
          6606 => x"ff",
          6607 => x"80",
          6608 => x"c0",
          6609 => x"87",
          6610 => x"bf",
          6611 => x"74",
          6612 => x"06",
          6613 => x"27",
          6614 => x"14",
          6615 => x"34",
          6616 => x"18",
          6617 => x"57",
          6618 => x"e3",
          6619 => x"ec",
          6620 => x"80",
          6621 => x"80",
          6622 => x"38",
          6623 => x"73",
          6624 => x"38",
          6625 => x"33",
          6626 => x"e0",
          6627 => x"d8",
          6628 => x"8c",
          6629 => x"54",
          6630 => x"94",
          6631 => x"55",
          6632 => x"74",
          6633 => x"38",
          6634 => x"33",
          6635 => x"39",
          6636 => x"05",
          6637 => x"78",
          6638 => x"56",
          6639 => x"76",
          6640 => x"38",
          6641 => x"15",
          6642 => x"55",
          6643 => x"34",
          6644 => x"e3",
          6645 => x"f9",
          6646 => x"d6",
          6647 => x"38",
          6648 => x"80",
          6649 => x"fe",
          6650 => x"55",
          6651 => x"2e",
          6652 => x"82",
          6653 => x"55",
          6654 => x"08",
          6655 => x"81",
          6656 => x"38",
          6657 => x"05",
          6658 => x"34",
          6659 => x"05",
          6660 => x"2a",
          6661 => x"51",
          6662 => x"59",
          6663 => x"90",
          6664 => x"8c",
          6665 => x"f8",
          6666 => x"d6",
          6667 => x"59",
          6668 => x"51",
          6669 => x"82",
          6670 => x"57",
          6671 => x"08",
          6672 => x"ff",
          6673 => x"80",
          6674 => x"38",
          6675 => x"90",
          6676 => x"31",
          6677 => x"51",
          6678 => x"82",
          6679 => x"57",
          6680 => x"08",
          6681 => x"a0",
          6682 => x"91",
          6683 => x"d8",
          6684 => x"06",
          6685 => x"08",
          6686 => x"e3",
          6687 => x"d6",
          6688 => x"82",
          6689 => x"81",
          6690 => x"1c",
          6691 => x"08",
          6692 => x"06",
          6693 => x"7c",
          6694 => x"8f",
          6695 => x"34",
          6696 => x"08",
          6697 => x"82",
          6698 => x"52",
          6699 => x"df",
          6700 => x"8d",
          6701 => x"77",
          6702 => x"83",
          6703 => x"8b",
          6704 => x"1b",
          6705 => x"17",
          6706 => x"73",
          6707 => x"d4",
          6708 => x"05",
          6709 => x"3f",
          6710 => x"83",
          6711 => x"81",
          6712 => x"77",
          6713 => x"73",
          6714 => x"2e",
          6715 => x"10",
          6716 => x"51",
          6717 => x"38",
          6718 => x"07",
          6719 => x"34",
          6720 => x"1d",
          6721 => x"79",
          6722 => x"3f",
          6723 => x"08",
          6724 => x"d8",
          6725 => x"38",
          6726 => x"78",
          6727 => x"98",
          6728 => x"7b",
          6729 => x"3f",
          6730 => x"08",
          6731 => x"d8",
          6732 => x"a0",
          6733 => x"d8",
          6734 => x"1a",
          6735 => x"c0",
          6736 => x"a0",
          6737 => x"1a",
          6738 => x"91",
          6739 => x"08",
          6740 => x"98",
          6741 => x"73",
          6742 => x"81",
          6743 => x"34",
          6744 => x"82",
          6745 => x"94",
          6746 => x"fa",
          6747 => x"70",
          6748 => x"08",
          6749 => x"56",
          6750 => x"72",
          6751 => x"38",
          6752 => x"51",
          6753 => x"82",
          6754 => x"54",
          6755 => x"08",
          6756 => x"98",
          6757 => x"75",
          6758 => x"3f",
          6759 => x"08",
          6760 => x"d8",
          6761 => x"9c",
          6762 => x"e5",
          6763 => x"0b",
          6764 => x"90",
          6765 => x"27",
          6766 => x"d6",
          6767 => x"74",
          6768 => x"3f",
          6769 => x"08",
          6770 => x"d8",
          6771 => x"c3",
          6772 => x"2e",
          6773 => x"83",
          6774 => x"73",
          6775 => x"0c",
          6776 => x"04",
          6777 => x"7e",
          6778 => x"5f",
          6779 => x"0b",
          6780 => x"98",
          6781 => x"2e",
          6782 => x"ac",
          6783 => x"2e",
          6784 => x"80",
          6785 => x"8c",
          6786 => x"22",
          6787 => x"5c",
          6788 => x"2e",
          6789 => x"78",
          6790 => x"22",
          6791 => x"56",
          6792 => x"38",
          6793 => x"15",
          6794 => x"ff",
          6795 => x"72",
          6796 => x"86",
          6797 => x"80",
          6798 => x"18",
          6799 => x"ff",
          6800 => x"5b",
          6801 => x"52",
          6802 => x"75",
          6803 => x"d5",
          6804 => x"d6",
          6805 => x"ff",
          6806 => x"81",
          6807 => x"95",
          6808 => x"27",
          6809 => x"88",
          6810 => x"7a",
          6811 => x"15",
          6812 => x"9f",
          6813 => x"76",
          6814 => x"07",
          6815 => x"80",
          6816 => x"54",
          6817 => x"2e",
          6818 => x"57",
          6819 => x"7a",
          6820 => x"74",
          6821 => x"5b",
          6822 => x"79",
          6823 => x"22",
          6824 => x"72",
          6825 => x"7a",
          6826 => x"25",
          6827 => x"06",
          6828 => x"77",
          6829 => x"53",
          6830 => x"14",
          6831 => x"89",
          6832 => x"57",
          6833 => x"19",
          6834 => x"1b",
          6835 => x"74",
          6836 => x"38",
          6837 => x"09",
          6838 => x"38",
          6839 => x"78",
          6840 => x"30",
          6841 => x"80",
          6842 => x"54",
          6843 => x"90",
          6844 => x"2e",
          6845 => x"76",
          6846 => x"58",
          6847 => x"57",
          6848 => x"81",
          6849 => x"81",
          6850 => x"79",
          6851 => x"38",
          6852 => x"05",
          6853 => x"81",
          6854 => x"18",
          6855 => x"81",
          6856 => x"8b",
          6857 => x"96",
          6858 => x"57",
          6859 => x"72",
          6860 => x"33",
          6861 => x"72",
          6862 => x"d3",
          6863 => x"89",
          6864 => x"73",
          6865 => x"11",
          6866 => x"99",
          6867 => x"9c",
          6868 => x"11",
          6869 => x"88",
          6870 => x"38",
          6871 => x"53",
          6872 => x"83",
          6873 => x"81",
          6874 => x"80",
          6875 => x"a0",
          6876 => x"ff",
          6877 => x"53",
          6878 => x"81",
          6879 => x"81",
          6880 => x"81",
          6881 => x"56",
          6882 => x"72",
          6883 => x"77",
          6884 => x"53",
          6885 => x"14",
          6886 => x"08",
          6887 => x"51",
          6888 => x"38",
          6889 => x"34",
          6890 => x"53",
          6891 => x"88",
          6892 => x"1c",
          6893 => x"52",
          6894 => x"3f",
          6895 => x"08",
          6896 => x"13",
          6897 => x"3f",
          6898 => x"08",
          6899 => x"98",
          6900 => x"fa",
          6901 => x"d8",
          6902 => x"23",
          6903 => x"04",
          6904 => x"62",
          6905 => x"5e",
          6906 => x"33",
          6907 => x"73",
          6908 => x"38",
          6909 => x"80",
          6910 => x"38",
          6911 => x"8d",
          6912 => x"05",
          6913 => x"0c",
          6914 => x"15",
          6915 => x"70",
          6916 => x"56",
          6917 => x"09",
          6918 => x"38",
          6919 => x"80",
          6920 => x"30",
          6921 => x"78",
          6922 => x"54",
          6923 => x"73",
          6924 => x"63",
          6925 => x"54",
          6926 => x"96",
          6927 => x"0b",
          6928 => x"80",
          6929 => x"e7",
          6930 => x"d6",
          6931 => x"87",
          6932 => x"41",
          6933 => x"11",
          6934 => x"80",
          6935 => x"fc",
          6936 => x"8f",
          6937 => x"d8",
          6938 => x"82",
          6939 => x"ff",
          6940 => x"d6",
          6941 => x"92",
          6942 => x"1a",
          6943 => x"08",
          6944 => x"55",
          6945 => x"81",
          6946 => x"d6",
          6947 => x"ff",
          6948 => x"af",
          6949 => x"9f",
          6950 => x"80",
          6951 => x"51",
          6952 => x"b4",
          6953 => x"dc",
          6954 => x"75",
          6955 => x"91",
          6956 => x"82",
          6957 => x"d9",
          6958 => x"d6",
          6959 => x"de",
          6960 => x"fe",
          6961 => x"38",
          6962 => x"54",
          6963 => x"81",
          6964 => x"89",
          6965 => x"41",
          6966 => x"33",
          6967 => x"73",
          6968 => x"81",
          6969 => x"81",
          6970 => x"dc",
          6971 => x"70",
          6972 => x"07",
          6973 => x"73",
          6974 => x"44",
          6975 => x"82",
          6976 => x"81",
          6977 => x"06",
          6978 => x"22",
          6979 => x"2e",
          6980 => x"d2",
          6981 => x"2e",
          6982 => x"80",
          6983 => x"1a",
          6984 => x"ae",
          6985 => x"06",
          6986 => x"79",
          6987 => x"ae",
          6988 => x"06",
          6989 => x"10",
          6990 => x"74",
          6991 => x"a0",
          6992 => x"ae",
          6993 => x"26",
          6994 => x"54",
          6995 => x"81",
          6996 => x"81",
          6997 => x"78",
          6998 => x"76",
          6999 => x"73",
          7000 => x"84",
          7001 => x"80",
          7002 => x"78",
          7003 => x"05",
          7004 => x"fe",
          7005 => x"a0",
          7006 => x"70",
          7007 => x"51",
          7008 => x"54",
          7009 => x"84",
          7010 => x"38",
          7011 => x"78",
          7012 => x"19",
          7013 => x"56",
          7014 => x"78",
          7015 => x"56",
          7016 => x"76",
          7017 => x"83",
          7018 => x"7a",
          7019 => x"ff",
          7020 => x"56",
          7021 => x"2e",
          7022 => x"93",
          7023 => x"70",
          7024 => x"22",
          7025 => x"73",
          7026 => x"38",
          7027 => x"74",
          7028 => x"06",
          7029 => x"2e",
          7030 => x"85",
          7031 => x"07",
          7032 => x"2e",
          7033 => x"16",
          7034 => x"22",
          7035 => x"ae",
          7036 => x"78",
          7037 => x"05",
          7038 => x"59",
          7039 => x"8f",
          7040 => x"70",
          7041 => x"73",
          7042 => x"81",
          7043 => x"8b",
          7044 => x"a0",
          7045 => x"e8",
          7046 => x"59",
          7047 => x"7c",
          7048 => x"22",
          7049 => x"57",
          7050 => x"2e",
          7051 => x"75",
          7052 => x"38",
          7053 => x"70",
          7054 => x"25",
          7055 => x"7c",
          7056 => x"38",
          7057 => x"89",
          7058 => x"07",
          7059 => x"80",
          7060 => x"7e",
          7061 => x"38",
          7062 => x"79",
          7063 => x"70",
          7064 => x"25",
          7065 => x"51",
          7066 => x"73",
          7067 => x"38",
          7068 => x"fe",
          7069 => x"79",
          7070 => x"76",
          7071 => x"7c",
          7072 => x"be",
          7073 => x"88",
          7074 => x"82",
          7075 => x"06",
          7076 => x"8b",
          7077 => x"76",
          7078 => x"76",
          7079 => x"83",
          7080 => x"51",
          7081 => x"3f",
          7082 => x"08",
          7083 => x"06",
          7084 => x"70",
          7085 => x"55",
          7086 => x"2e",
          7087 => x"80",
          7088 => x"c7",
          7089 => x"57",
          7090 => x"76",
          7091 => x"ff",
          7092 => x"78",
          7093 => x"76",
          7094 => x"59",
          7095 => x"39",
          7096 => x"05",
          7097 => x"55",
          7098 => x"34",
          7099 => x"80",
          7100 => x"80",
          7101 => x"75",
          7102 => x"fc",
          7103 => x"3f",
          7104 => x"08",
          7105 => x"38",
          7106 => x"83",
          7107 => x"a4",
          7108 => x"16",
          7109 => x"26",
          7110 => x"82",
          7111 => x"9f",
          7112 => x"99",
          7113 => x"7b",
          7114 => x"17",
          7115 => x"ff",
          7116 => x"5c",
          7117 => x"05",
          7118 => x"34",
          7119 => x"fd",
          7120 => x"1e",
          7121 => x"81",
          7122 => x"81",
          7123 => x"85",
          7124 => x"34",
          7125 => x"09",
          7126 => x"38",
          7127 => x"81",
          7128 => x"7b",
          7129 => x"73",
          7130 => x"38",
          7131 => x"54",
          7132 => x"09",
          7133 => x"38",
          7134 => x"57",
          7135 => x"70",
          7136 => x"54",
          7137 => x"7b",
          7138 => x"73",
          7139 => x"38",
          7140 => x"57",
          7141 => x"70",
          7142 => x"54",
          7143 => x"85",
          7144 => x"07",
          7145 => x"1f",
          7146 => x"ea",
          7147 => x"d6",
          7148 => x"1f",
          7149 => x"82",
          7150 => x"80",
          7151 => x"82",
          7152 => x"84",
          7153 => x"06",
          7154 => x"74",
          7155 => x"81",
          7156 => x"2a",
          7157 => x"73",
          7158 => x"38",
          7159 => x"54",
          7160 => x"f8",
          7161 => x"80",
          7162 => x"34",
          7163 => x"c2",
          7164 => x"06",
          7165 => x"38",
          7166 => x"39",
          7167 => x"70",
          7168 => x"54",
          7169 => x"86",
          7170 => x"84",
          7171 => x"06",
          7172 => x"73",
          7173 => x"38",
          7174 => x"83",
          7175 => x"05",
          7176 => x"7f",
          7177 => x"3f",
          7178 => x"08",
          7179 => x"f8",
          7180 => x"82",
          7181 => x"92",
          7182 => x"f6",
          7183 => x"5b",
          7184 => x"70",
          7185 => x"59",
          7186 => x"73",
          7187 => x"c6",
          7188 => x"81",
          7189 => x"70",
          7190 => x"52",
          7191 => x"8d",
          7192 => x"38",
          7193 => x"09",
          7194 => x"a5",
          7195 => x"d0",
          7196 => x"ff",
          7197 => x"53",
          7198 => x"91",
          7199 => x"73",
          7200 => x"d0",
          7201 => x"71",
          7202 => x"f7",
          7203 => x"82",
          7204 => x"55",
          7205 => x"55",
          7206 => x"81",
          7207 => x"74",
          7208 => x"56",
          7209 => x"12",
          7210 => x"70",
          7211 => x"38",
          7212 => x"81",
          7213 => x"51",
          7214 => x"51",
          7215 => x"89",
          7216 => x"70",
          7217 => x"53",
          7218 => x"70",
          7219 => x"51",
          7220 => x"09",
          7221 => x"38",
          7222 => x"38",
          7223 => x"77",
          7224 => x"70",
          7225 => x"2a",
          7226 => x"07",
          7227 => x"51",
          7228 => x"8f",
          7229 => x"84",
          7230 => x"83",
          7231 => x"94",
          7232 => x"74",
          7233 => x"38",
          7234 => x"0c",
          7235 => x"86",
          7236 => x"b4",
          7237 => x"82",
          7238 => x"8c",
          7239 => x"fa",
          7240 => x"56",
          7241 => x"17",
          7242 => x"b4",
          7243 => x"52",
          7244 => x"f4",
          7245 => x"82",
          7246 => x"81",
          7247 => x"b6",
          7248 => x"8a",
          7249 => x"d8",
          7250 => x"ff",
          7251 => x"55",
          7252 => x"d5",
          7253 => x"06",
          7254 => x"80",
          7255 => x"33",
          7256 => x"81",
          7257 => x"81",
          7258 => x"81",
          7259 => x"eb",
          7260 => x"70",
          7261 => x"07",
          7262 => x"73",
          7263 => x"81",
          7264 => x"81",
          7265 => x"83",
          7266 => x"84",
          7267 => x"16",
          7268 => x"3f",
          7269 => x"08",
          7270 => x"d8",
          7271 => x"9d",
          7272 => x"82",
          7273 => x"81",
          7274 => x"ce",
          7275 => x"d6",
          7276 => x"82",
          7277 => x"80",
          7278 => x"82",
          7279 => x"d6",
          7280 => x"3d",
          7281 => x"3d",
          7282 => x"84",
          7283 => x"05",
          7284 => x"80",
          7285 => x"51",
          7286 => x"82",
          7287 => x"58",
          7288 => x"0b",
          7289 => x"08",
          7290 => x"38",
          7291 => x"08",
          7292 => x"ee",
          7293 => x"08",
          7294 => x"56",
          7295 => x"86",
          7296 => x"75",
          7297 => x"fe",
          7298 => x"54",
          7299 => x"2e",
          7300 => x"14",
          7301 => x"a0",
          7302 => x"d8",
          7303 => x"06",
          7304 => x"54",
          7305 => x"38",
          7306 => x"86",
          7307 => x"82",
          7308 => x"06",
          7309 => x"56",
          7310 => x"38",
          7311 => x"80",
          7312 => x"81",
          7313 => x"52",
          7314 => x"51",
          7315 => x"82",
          7316 => x"81",
          7317 => x"81",
          7318 => x"83",
          7319 => x"8f",
          7320 => x"2e",
          7321 => x"82",
          7322 => x"06",
          7323 => x"56",
          7324 => x"38",
          7325 => x"74",
          7326 => x"a3",
          7327 => x"d8",
          7328 => x"06",
          7329 => x"2e",
          7330 => x"80",
          7331 => x"3d",
          7332 => x"83",
          7333 => x"15",
          7334 => x"53",
          7335 => x"8d",
          7336 => x"15",
          7337 => x"3f",
          7338 => x"08",
          7339 => x"70",
          7340 => x"0c",
          7341 => x"16",
          7342 => x"80",
          7343 => x"80",
          7344 => x"54",
          7345 => x"84",
          7346 => x"5b",
          7347 => x"80",
          7348 => x"7a",
          7349 => x"fc",
          7350 => x"d6",
          7351 => x"ff",
          7352 => x"77",
          7353 => x"81",
          7354 => x"76",
          7355 => x"81",
          7356 => x"2e",
          7357 => x"8d",
          7358 => x"26",
          7359 => x"80",
          7360 => x"ca",
          7361 => x"d6",
          7362 => x"ff",
          7363 => x"72",
          7364 => x"09",
          7365 => x"d7",
          7366 => x"14",
          7367 => x"3f",
          7368 => x"08",
          7369 => x"06",
          7370 => x"38",
          7371 => x"51",
          7372 => x"82",
          7373 => x"58",
          7374 => x"0c",
          7375 => x"33",
          7376 => x"80",
          7377 => x"ff",
          7378 => x"ff",
          7379 => x"55",
          7380 => x"81",
          7381 => x"38",
          7382 => x"06",
          7383 => x"80",
          7384 => x"52",
          7385 => x"8a",
          7386 => x"80",
          7387 => x"ff",
          7388 => x"53",
          7389 => x"86",
          7390 => x"83",
          7391 => x"c9",
          7392 => x"ca",
          7393 => x"d8",
          7394 => x"d6",
          7395 => x"15",
          7396 => x"06",
          7397 => x"76",
          7398 => x"80",
          7399 => x"c9",
          7400 => x"d6",
          7401 => x"ff",
          7402 => x"74",
          7403 => x"d8",
          7404 => x"b1",
          7405 => x"d8",
          7406 => x"c6",
          7407 => x"8e",
          7408 => x"d8",
          7409 => x"ff",
          7410 => x"56",
          7411 => x"83",
          7412 => x"14",
          7413 => x"71",
          7414 => x"5a",
          7415 => x"26",
          7416 => x"8a",
          7417 => x"74",
          7418 => x"fe",
          7419 => x"82",
          7420 => x"55",
          7421 => x"08",
          7422 => x"f3",
          7423 => x"d8",
          7424 => x"ff",
          7425 => x"83",
          7426 => x"74",
          7427 => x"26",
          7428 => x"57",
          7429 => x"26",
          7430 => x"57",
          7431 => x"56",
          7432 => x"82",
          7433 => x"15",
          7434 => x"0c",
          7435 => x"0c",
          7436 => x"a8",
          7437 => x"1d",
          7438 => x"54",
          7439 => x"2e",
          7440 => x"af",
          7441 => x"14",
          7442 => x"3f",
          7443 => x"08",
          7444 => x"06",
          7445 => x"72",
          7446 => x"79",
          7447 => x"80",
          7448 => x"c8",
          7449 => x"d6",
          7450 => x"15",
          7451 => x"2b",
          7452 => x"8d",
          7453 => x"2e",
          7454 => x"77",
          7455 => x"0c",
          7456 => x"76",
          7457 => x"38",
          7458 => x"70",
          7459 => x"81",
          7460 => x"53",
          7461 => x"89",
          7462 => x"56",
          7463 => x"08",
          7464 => x"38",
          7465 => x"15",
          7466 => x"90",
          7467 => x"80",
          7468 => x"34",
          7469 => x"09",
          7470 => x"92",
          7471 => x"14",
          7472 => x"3f",
          7473 => x"08",
          7474 => x"06",
          7475 => x"2e",
          7476 => x"80",
          7477 => x"1b",
          7478 => x"ca",
          7479 => x"d6",
          7480 => x"ea",
          7481 => x"d8",
          7482 => x"34",
          7483 => x"51",
          7484 => x"82",
          7485 => x"83",
          7486 => x"53",
          7487 => x"d5",
          7488 => x"06",
          7489 => x"b8",
          7490 => x"d9",
          7491 => x"d8",
          7492 => x"85",
          7493 => x"09",
          7494 => x"38",
          7495 => x"51",
          7496 => x"82",
          7497 => x"86",
          7498 => x"f2",
          7499 => x"06",
          7500 => x"a0",
          7501 => x"ad",
          7502 => x"d8",
          7503 => x"0c",
          7504 => x"51",
          7505 => x"82",
          7506 => x"90",
          7507 => x"74",
          7508 => x"b0",
          7509 => x"53",
          7510 => x"b0",
          7511 => x"15",
          7512 => x"b8",
          7513 => x"0c",
          7514 => x"15",
          7515 => x"75",
          7516 => x"0c",
          7517 => x"04",
          7518 => x"77",
          7519 => x"73",
          7520 => x"38",
          7521 => x"72",
          7522 => x"38",
          7523 => x"71",
          7524 => x"38",
          7525 => x"84",
          7526 => x"52",
          7527 => x"09",
          7528 => x"38",
          7529 => x"51",
          7530 => x"3f",
          7531 => x"08",
          7532 => x"71",
          7533 => x"74",
          7534 => x"83",
          7535 => x"78",
          7536 => x"52",
          7537 => x"d8",
          7538 => x"0d",
          7539 => x"0d",
          7540 => x"33",
          7541 => x"3d",
          7542 => x"56",
          7543 => x"8b",
          7544 => x"82",
          7545 => x"24",
          7546 => x"d6",
          7547 => x"29",
          7548 => x"05",
          7549 => x"55",
          7550 => x"84",
          7551 => x"34",
          7552 => x"80",
          7553 => x"80",
          7554 => x"75",
          7555 => x"75",
          7556 => x"38",
          7557 => x"3d",
          7558 => x"05",
          7559 => x"3f",
          7560 => x"08",
          7561 => x"d6",
          7562 => x"3d",
          7563 => x"3d",
          7564 => x"84",
          7565 => x"05",
          7566 => x"89",
          7567 => x"2e",
          7568 => x"77",
          7569 => x"54",
          7570 => x"05",
          7571 => x"84",
          7572 => x"f6",
          7573 => x"d6",
          7574 => x"82",
          7575 => x"84",
          7576 => x"5c",
          7577 => x"3d",
          7578 => x"ea",
          7579 => x"d6",
          7580 => x"82",
          7581 => x"92",
          7582 => x"d7",
          7583 => x"98",
          7584 => x"73",
          7585 => x"38",
          7586 => x"9c",
          7587 => x"80",
          7588 => x"38",
          7589 => x"95",
          7590 => x"2e",
          7591 => x"aa",
          7592 => x"df",
          7593 => x"d6",
          7594 => x"9e",
          7595 => x"05",
          7596 => x"54",
          7597 => x"38",
          7598 => x"70",
          7599 => x"54",
          7600 => x"8e",
          7601 => x"83",
          7602 => x"88",
          7603 => x"83",
          7604 => x"83",
          7605 => x"06",
          7606 => x"80",
          7607 => x"38",
          7608 => x"51",
          7609 => x"82",
          7610 => x"56",
          7611 => x"0a",
          7612 => x"05",
          7613 => x"3f",
          7614 => x"0b",
          7615 => x"80",
          7616 => x"7a",
          7617 => x"3f",
          7618 => x"9c",
          7619 => x"9e",
          7620 => x"81",
          7621 => x"34",
          7622 => x"80",
          7623 => x"b4",
          7624 => x"54",
          7625 => x"52",
          7626 => x"05",
          7627 => x"3f",
          7628 => x"08",
          7629 => x"d8",
          7630 => x"38",
          7631 => x"82",
          7632 => x"b2",
          7633 => x"84",
          7634 => x"06",
          7635 => x"73",
          7636 => x"38",
          7637 => x"ad",
          7638 => x"2a",
          7639 => x"51",
          7640 => x"2e",
          7641 => x"81",
          7642 => x"80",
          7643 => x"87",
          7644 => x"39",
          7645 => x"51",
          7646 => x"82",
          7647 => x"7b",
          7648 => x"12",
          7649 => x"82",
          7650 => x"81",
          7651 => x"83",
          7652 => x"06",
          7653 => x"80",
          7654 => x"77",
          7655 => x"58",
          7656 => x"08",
          7657 => x"63",
          7658 => x"63",
          7659 => x"57",
          7660 => x"82",
          7661 => x"82",
          7662 => x"88",
          7663 => x"9c",
          7664 => x"c1",
          7665 => x"d6",
          7666 => x"d6",
          7667 => x"1b",
          7668 => x"0c",
          7669 => x"22",
          7670 => x"77",
          7671 => x"80",
          7672 => x"34",
          7673 => x"1a",
          7674 => x"94",
          7675 => x"85",
          7676 => x"06",
          7677 => x"80",
          7678 => x"38",
          7679 => x"08",
          7680 => x"84",
          7681 => x"d8",
          7682 => x"0c",
          7683 => x"70",
          7684 => x"52",
          7685 => x"39",
          7686 => x"51",
          7687 => x"82",
          7688 => x"57",
          7689 => x"08",
          7690 => x"38",
          7691 => x"d6",
          7692 => x"2e",
          7693 => x"83",
          7694 => x"75",
          7695 => x"74",
          7696 => x"07",
          7697 => x"54",
          7698 => x"8a",
          7699 => x"75",
          7700 => x"73",
          7701 => x"98",
          7702 => x"a9",
          7703 => x"ff",
          7704 => x"80",
          7705 => x"76",
          7706 => x"c5",
          7707 => x"d6",
          7708 => x"38",
          7709 => x"39",
          7710 => x"82",
          7711 => x"05",
          7712 => x"84",
          7713 => x"0c",
          7714 => x"82",
          7715 => x"98",
          7716 => x"f2",
          7717 => x"63",
          7718 => x"40",
          7719 => x"7e",
          7720 => x"fc",
          7721 => x"51",
          7722 => x"82",
          7723 => x"55",
          7724 => x"08",
          7725 => x"19",
          7726 => x"80",
          7727 => x"74",
          7728 => x"39",
          7729 => x"81",
          7730 => x"56",
          7731 => x"82",
          7732 => x"39",
          7733 => x"1a",
          7734 => x"82",
          7735 => x"0b",
          7736 => x"81",
          7737 => x"39",
          7738 => x"94",
          7739 => x"55",
          7740 => x"83",
          7741 => x"7b",
          7742 => x"8c",
          7743 => x"08",
          7744 => x"06",
          7745 => x"81",
          7746 => x"8a",
          7747 => x"05",
          7748 => x"06",
          7749 => x"a8",
          7750 => x"38",
          7751 => x"55",
          7752 => x"19",
          7753 => x"51",
          7754 => x"82",
          7755 => x"55",
          7756 => x"ff",
          7757 => x"ff",
          7758 => x"38",
          7759 => x"0c",
          7760 => x"52",
          7761 => x"d6",
          7762 => x"d8",
          7763 => x"ff",
          7764 => x"d6",
          7765 => x"7c",
          7766 => x"57",
          7767 => x"80",
          7768 => x"1a",
          7769 => x"22",
          7770 => x"75",
          7771 => x"38",
          7772 => x"58",
          7773 => x"53",
          7774 => x"1b",
          7775 => x"b8",
          7776 => x"d6",
          7777 => x"d6",
          7778 => x"11",
          7779 => x"74",
          7780 => x"38",
          7781 => x"77",
          7782 => x"78",
          7783 => x"84",
          7784 => x"16",
          7785 => x"08",
          7786 => x"2b",
          7787 => x"ff",
          7788 => x"77",
          7789 => x"ba",
          7790 => x"1a",
          7791 => x"08",
          7792 => x"84",
          7793 => x"57",
          7794 => x"27",
          7795 => x"56",
          7796 => x"52",
          7797 => x"d0",
          7798 => x"d8",
          7799 => x"38",
          7800 => x"19",
          7801 => x"06",
          7802 => x"52",
          7803 => x"bd",
          7804 => x"76",
          7805 => x"17",
          7806 => x"1e",
          7807 => x"18",
          7808 => x"5e",
          7809 => x"39",
          7810 => x"82",
          7811 => x"90",
          7812 => x"f2",
          7813 => x"63",
          7814 => x"40",
          7815 => x"7e",
          7816 => x"fc",
          7817 => x"51",
          7818 => x"82",
          7819 => x"55",
          7820 => x"08",
          7821 => x"18",
          7822 => x"80",
          7823 => x"74",
          7824 => x"39",
          7825 => x"70",
          7826 => x"81",
          7827 => x"56",
          7828 => x"80",
          7829 => x"38",
          7830 => x"0b",
          7831 => x"82",
          7832 => x"39",
          7833 => x"19",
          7834 => x"83",
          7835 => x"18",
          7836 => x"56",
          7837 => x"27",
          7838 => x"09",
          7839 => x"2e",
          7840 => x"94",
          7841 => x"83",
          7842 => x"56",
          7843 => x"38",
          7844 => x"22",
          7845 => x"89",
          7846 => x"55",
          7847 => x"75",
          7848 => x"18",
          7849 => x"9c",
          7850 => x"85",
          7851 => x"08",
          7852 => x"c6",
          7853 => x"d6",
          7854 => x"82",
          7855 => x"80",
          7856 => x"38",
          7857 => x"ff",
          7858 => x"ff",
          7859 => x"38",
          7860 => x"0c",
          7861 => x"85",
          7862 => x"19",
          7863 => x"b4",
          7864 => x"19",
          7865 => x"81",
          7866 => x"74",
          7867 => x"c8",
          7868 => x"d8",
          7869 => x"38",
          7870 => x"52",
          7871 => x"9e",
          7872 => x"d8",
          7873 => x"fe",
          7874 => x"d6",
          7875 => x"7c",
          7876 => x"57",
          7877 => x"80",
          7878 => x"1b",
          7879 => x"22",
          7880 => x"75",
          7881 => x"38",
          7882 => x"59",
          7883 => x"53",
          7884 => x"1a",
          7885 => x"b7",
          7886 => x"d6",
          7887 => x"a4",
          7888 => x"11",
          7889 => x"56",
          7890 => x"27",
          7891 => x"80",
          7892 => x"08",
          7893 => x"2b",
          7894 => x"b8",
          7895 => x"ba",
          7896 => x"55",
          7897 => x"16",
          7898 => x"2b",
          7899 => x"39",
          7900 => x"94",
          7901 => x"94",
          7902 => x"ff",
          7903 => x"82",
          7904 => x"fd",
          7905 => x"77",
          7906 => x"55",
          7907 => x"0c",
          7908 => x"83",
          7909 => x"80",
          7910 => x"55",
          7911 => x"83",
          7912 => x"9c",
          7913 => x"7e",
          7914 => x"fc",
          7915 => x"d8",
          7916 => x"38",
          7917 => x"52",
          7918 => x"83",
          7919 => x"b8",
          7920 => x"ba",
          7921 => x"55",
          7922 => x"16",
          7923 => x"31",
          7924 => x"7f",
          7925 => x"94",
          7926 => x"70",
          7927 => x"8c",
          7928 => x"58",
          7929 => x"76",
          7930 => x"75",
          7931 => x"19",
          7932 => x"39",
          7933 => x"80",
          7934 => x"74",
          7935 => x"80",
          7936 => x"d6",
          7937 => x"3d",
          7938 => x"3d",
          7939 => x"3d",
          7940 => x"70",
          7941 => x"e0",
          7942 => x"d8",
          7943 => x"d6",
          7944 => x"80",
          7945 => x"33",
          7946 => x"70",
          7947 => x"55",
          7948 => x"2e",
          7949 => x"a0",
          7950 => x"78",
          7951 => x"e8",
          7952 => x"d8",
          7953 => x"d6",
          7954 => x"d8",
          7955 => x"08",
          7956 => x"a0",
          7957 => x"73",
          7958 => x"88",
          7959 => x"74",
          7960 => x"51",
          7961 => x"8c",
          7962 => x"9c",
          7963 => x"b8",
          7964 => x"88",
          7965 => x"96",
          7966 => x"b8",
          7967 => x"52",
          7968 => x"ff",
          7969 => x"78",
          7970 => x"83",
          7971 => x"51",
          7972 => x"3f",
          7973 => x"08",
          7974 => x"81",
          7975 => x"57",
          7976 => x"34",
          7977 => x"d8",
          7978 => x"0d",
          7979 => x"0d",
          7980 => x"54",
          7981 => x"82",
          7982 => x"53",
          7983 => x"08",
          7984 => x"3d",
          7985 => x"73",
          7986 => x"3f",
          7987 => x"08",
          7988 => x"d8",
          7989 => x"82",
          7990 => x"74",
          7991 => x"d6",
          7992 => x"3d",
          7993 => x"3d",
          7994 => x"51",
          7995 => x"8b",
          7996 => x"82",
          7997 => x"24",
          7998 => x"d6",
          7999 => x"ee",
          8000 => x"52",
          8001 => x"d8",
          8002 => x"0d",
          8003 => x"0d",
          8004 => x"3d",
          8005 => x"95",
          8006 => x"aa",
          8007 => x"d8",
          8008 => x"d6",
          8009 => x"e0",
          8010 => x"64",
          8011 => x"d0",
          8012 => x"ac",
          8013 => x"d8",
          8014 => x"d6",
          8015 => x"38",
          8016 => x"05",
          8017 => x"2b",
          8018 => x"80",
          8019 => x"76",
          8020 => x"0c",
          8021 => x"02",
          8022 => x"70",
          8023 => x"81",
          8024 => x"56",
          8025 => x"9e",
          8026 => x"53",
          8027 => x"ca",
          8028 => x"d6",
          8029 => x"15",
          8030 => x"82",
          8031 => x"84",
          8032 => x"06",
          8033 => x"55",
          8034 => x"d8",
          8035 => x"0d",
          8036 => x"3d",
          8037 => x"3d",
          8038 => x"3d",
          8039 => x"80",
          8040 => x"53",
          8041 => x"fd",
          8042 => x"80",
          8043 => x"e8",
          8044 => x"d6",
          8045 => x"82",
          8046 => x"83",
          8047 => x"80",
          8048 => x"7a",
          8049 => x"08",
          8050 => x"0c",
          8051 => x"d5",
          8052 => x"73",
          8053 => x"83",
          8054 => x"80",
          8055 => x"52",
          8056 => x"3f",
          8057 => x"08",
          8058 => x"d8",
          8059 => x"38",
          8060 => x"08",
          8061 => x"ff",
          8062 => x"82",
          8063 => x"57",
          8064 => x"08",
          8065 => x"80",
          8066 => x"52",
          8067 => x"86",
          8068 => x"d8",
          8069 => x"3d",
          8070 => x"74",
          8071 => x"3f",
          8072 => x"08",
          8073 => x"d8",
          8074 => x"38",
          8075 => x"51",
          8076 => x"82",
          8077 => x"57",
          8078 => x"08",
          8079 => x"da",
          8080 => x"7b",
          8081 => x"3f",
          8082 => x"d8",
          8083 => x"38",
          8084 => x"51",
          8085 => x"82",
          8086 => x"57",
          8087 => x"08",
          8088 => x"38",
          8089 => x"09",
          8090 => x"38",
          8091 => x"ee",
          8092 => x"ea",
          8093 => x"3d",
          8094 => x"52",
          8095 => x"e4",
          8096 => x"3d",
          8097 => x"11",
          8098 => x"5a",
          8099 => x"2e",
          8100 => x"80",
          8101 => x"81",
          8102 => x"70",
          8103 => x"56",
          8104 => x"81",
          8105 => x"78",
          8106 => x"38",
          8107 => x"9c",
          8108 => x"82",
          8109 => x"18",
          8110 => x"08",
          8111 => x"ff",
          8112 => x"55",
          8113 => x"74",
          8114 => x"38",
          8115 => x"e1",
          8116 => x"55",
          8117 => x"34",
          8118 => x"77",
          8119 => x"81",
          8120 => x"ff",
          8121 => x"3d",
          8122 => x"58",
          8123 => x"80",
          8124 => x"b4",
          8125 => x"29",
          8126 => x"05",
          8127 => x"33",
          8128 => x"56",
          8129 => x"2e",
          8130 => x"16",
          8131 => x"33",
          8132 => x"73",
          8133 => x"16",
          8134 => x"26",
          8135 => x"55",
          8136 => x"91",
          8137 => x"54",
          8138 => x"70",
          8139 => x"34",
          8140 => x"ec",
          8141 => x"70",
          8142 => x"34",
          8143 => x"09",
          8144 => x"38",
          8145 => x"39",
          8146 => x"08",
          8147 => x"59",
          8148 => x"7a",
          8149 => x"5c",
          8150 => x"26",
          8151 => x"7a",
          8152 => x"d6",
          8153 => x"df",
          8154 => x"f7",
          8155 => x"7d",
          8156 => x"05",
          8157 => x"57",
          8158 => x"3f",
          8159 => x"08",
          8160 => x"d8",
          8161 => x"38",
          8162 => x"53",
          8163 => x"38",
          8164 => x"54",
          8165 => x"92",
          8166 => x"33",
          8167 => x"70",
          8168 => x"54",
          8169 => x"38",
          8170 => x"15",
          8171 => x"70",
          8172 => x"58",
          8173 => x"82",
          8174 => x"8a",
          8175 => x"89",
          8176 => x"53",
          8177 => x"b7",
          8178 => x"ff",
          8179 => x"c8",
          8180 => x"d6",
          8181 => x"15",
          8182 => x"53",
          8183 => x"c8",
          8184 => x"d6",
          8185 => x"26",
          8186 => x"30",
          8187 => x"70",
          8188 => x"77",
          8189 => x"18",
          8190 => x"51",
          8191 => x"88",
          8192 => x"73",
          8193 => x"52",
          8194 => x"bc",
          8195 => x"d6",
          8196 => x"82",
          8197 => x"81",
          8198 => x"38",
          8199 => x"08",
          8200 => x"9e",
          8201 => x"d8",
          8202 => x"0c",
          8203 => x"0c",
          8204 => x"81",
          8205 => x"76",
          8206 => x"38",
          8207 => x"94",
          8208 => x"94",
          8209 => x"16",
          8210 => x"2a",
          8211 => x"51",
          8212 => x"72",
          8213 => x"38",
          8214 => x"51",
          8215 => x"3f",
          8216 => x"08",
          8217 => x"d8",
          8218 => x"82",
          8219 => x"56",
          8220 => x"52",
          8221 => x"b5",
          8222 => x"d6",
          8223 => x"73",
          8224 => x"38",
          8225 => x"b0",
          8226 => x"73",
          8227 => x"27",
          8228 => x"98",
          8229 => x"9e",
          8230 => x"08",
          8231 => x"0c",
          8232 => x"06",
          8233 => x"2e",
          8234 => x"52",
          8235 => x"b4",
          8236 => x"d6",
          8237 => x"38",
          8238 => x"16",
          8239 => x"80",
          8240 => x"0b",
          8241 => x"81",
          8242 => x"75",
          8243 => x"d6",
          8244 => x"58",
          8245 => x"54",
          8246 => x"74",
          8247 => x"73",
          8248 => x"90",
          8249 => x"c0",
          8250 => x"90",
          8251 => x"83",
          8252 => x"72",
          8253 => x"38",
          8254 => x"08",
          8255 => x"77",
          8256 => x"80",
          8257 => x"d6",
          8258 => x"3d",
          8259 => x"3d",
          8260 => x"89",
          8261 => x"2e",
          8262 => x"80",
          8263 => x"fc",
          8264 => x"3d",
          8265 => x"e1",
          8266 => x"d6",
          8267 => x"82",
          8268 => x"80",
          8269 => x"76",
          8270 => x"75",
          8271 => x"3f",
          8272 => x"08",
          8273 => x"d8",
          8274 => x"38",
          8275 => x"70",
          8276 => x"57",
          8277 => x"a2",
          8278 => x"33",
          8279 => x"70",
          8280 => x"55",
          8281 => x"2e",
          8282 => x"16",
          8283 => x"51",
          8284 => x"82",
          8285 => x"88",
          8286 => x"54",
          8287 => x"84",
          8288 => x"52",
          8289 => x"bd",
          8290 => x"d6",
          8291 => x"74",
          8292 => x"81",
          8293 => x"85",
          8294 => x"74",
          8295 => x"38",
          8296 => x"74",
          8297 => x"d6",
          8298 => x"3d",
          8299 => x"3d",
          8300 => x"3d",
          8301 => x"70",
          8302 => x"bc",
          8303 => x"d8",
          8304 => x"82",
          8305 => x"73",
          8306 => x"0d",
          8307 => x"0d",
          8308 => x"3d",
          8309 => x"71",
          8310 => x"e7",
          8311 => x"d6",
          8312 => x"82",
          8313 => x"80",
          8314 => x"94",
          8315 => x"d8",
          8316 => x"51",
          8317 => x"3f",
          8318 => x"08",
          8319 => x"39",
          8320 => x"08",
          8321 => x"c2",
          8322 => x"d6",
          8323 => x"82",
          8324 => x"84",
          8325 => x"06",
          8326 => x"53",
          8327 => x"d6",
          8328 => x"38",
          8329 => x"51",
          8330 => x"72",
          8331 => x"ff",
          8332 => x"82",
          8333 => x"84",
          8334 => x"70",
          8335 => x"2c",
          8336 => x"d8",
          8337 => x"51",
          8338 => x"82",
          8339 => x"87",
          8340 => x"ed",
          8341 => x"57",
          8342 => x"3d",
          8343 => x"3d",
          8344 => x"e2",
          8345 => x"d8",
          8346 => x"d6",
          8347 => x"38",
          8348 => x"51",
          8349 => x"82",
          8350 => x"55",
          8351 => x"08",
          8352 => x"80",
          8353 => x"70",
          8354 => x"58",
          8355 => x"85",
          8356 => x"8d",
          8357 => x"2e",
          8358 => x"52",
          8359 => x"c4",
          8360 => x"d6",
          8361 => x"3d",
          8362 => x"3d",
          8363 => x"55",
          8364 => x"92",
          8365 => x"52",
          8366 => x"de",
          8367 => x"d6",
          8368 => x"82",
          8369 => x"82",
          8370 => x"74",
          8371 => x"9c",
          8372 => x"11",
          8373 => x"59",
          8374 => x"75",
          8375 => x"38",
          8376 => x"81",
          8377 => x"5b",
          8378 => x"82",
          8379 => x"39",
          8380 => x"08",
          8381 => x"59",
          8382 => x"09",
          8383 => x"c0",
          8384 => x"5f",
          8385 => x"92",
          8386 => x"51",
          8387 => x"3f",
          8388 => x"08",
          8389 => x"38",
          8390 => x"08",
          8391 => x"38",
          8392 => x"08",
          8393 => x"d6",
          8394 => x"80",
          8395 => x"81",
          8396 => x"59",
          8397 => x"14",
          8398 => x"c9",
          8399 => x"39",
          8400 => x"82",
          8401 => x"57",
          8402 => x"38",
          8403 => x"18",
          8404 => x"ff",
          8405 => x"82",
          8406 => x"5b",
          8407 => x"08",
          8408 => x"7c",
          8409 => x"12",
          8410 => x"52",
          8411 => x"82",
          8412 => x"06",
          8413 => x"14",
          8414 => x"d2",
          8415 => x"d8",
          8416 => x"ff",
          8417 => x"70",
          8418 => x"82",
          8419 => x"51",
          8420 => x"b8",
          8421 => x"a9",
          8422 => x"d6",
          8423 => x"0a",
          8424 => x"70",
          8425 => x"84",
          8426 => x"51",
          8427 => x"ff",
          8428 => x"56",
          8429 => x"38",
          8430 => x"7c",
          8431 => x"0c",
          8432 => x"81",
          8433 => x"74",
          8434 => x"7a",
          8435 => x"0c",
          8436 => x"04",
          8437 => x"79",
          8438 => x"05",
          8439 => x"57",
          8440 => x"82",
          8441 => x"56",
          8442 => x"08",
          8443 => x"91",
          8444 => x"75",
          8445 => x"90",
          8446 => x"81",
          8447 => x"06",
          8448 => x"87",
          8449 => x"2e",
          8450 => x"94",
          8451 => x"73",
          8452 => x"27",
          8453 => x"73",
          8454 => x"d6",
          8455 => x"88",
          8456 => x"76",
          8457 => x"d0",
          8458 => x"d8",
          8459 => x"19",
          8460 => x"ca",
          8461 => x"08",
          8462 => x"ff",
          8463 => x"82",
          8464 => x"ff",
          8465 => x"06",
          8466 => x"56",
          8467 => x"08",
          8468 => x"81",
          8469 => x"82",
          8470 => x"75",
          8471 => x"54",
          8472 => x"08",
          8473 => x"27",
          8474 => x"17",
          8475 => x"d6",
          8476 => x"76",
          8477 => x"80",
          8478 => x"d8",
          8479 => x"17",
          8480 => x"0c",
          8481 => x"80",
          8482 => x"73",
          8483 => x"75",
          8484 => x"38",
          8485 => x"34",
          8486 => x"82",
          8487 => x"89",
          8488 => x"e0",
          8489 => x"53",
          8490 => x"9c",
          8491 => x"3d",
          8492 => x"3f",
          8493 => x"08",
          8494 => x"d8",
          8495 => x"38",
          8496 => x"3d",
          8497 => x"3d",
          8498 => x"ce",
          8499 => x"d6",
          8500 => x"82",
          8501 => x"81",
          8502 => x"80",
          8503 => x"70",
          8504 => x"81",
          8505 => x"56",
          8506 => x"81",
          8507 => x"98",
          8508 => x"74",
          8509 => x"38",
          8510 => x"05",
          8511 => x"06",
          8512 => x"55",
          8513 => x"38",
          8514 => x"51",
          8515 => x"3f",
          8516 => x"08",
          8517 => x"70",
          8518 => x"55",
          8519 => x"2e",
          8520 => x"78",
          8521 => x"d8",
          8522 => x"08",
          8523 => x"38",
          8524 => x"d6",
          8525 => x"76",
          8526 => x"70",
          8527 => x"b5",
          8528 => x"d6",
          8529 => x"82",
          8530 => x"80",
          8531 => x"d6",
          8532 => x"73",
          8533 => x"d4",
          8534 => x"d8",
          8535 => x"d6",
          8536 => x"38",
          8537 => x"d0",
          8538 => x"d8",
          8539 => x"88",
          8540 => x"d8",
          8541 => x"38",
          8542 => x"ef",
          8543 => x"d8",
          8544 => x"d8",
          8545 => x"82",
          8546 => x"07",
          8547 => x"55",
          8548 => x"2e",
          8549 => x"80",
          8550 => x"80",
          8551 => x"77",
          8552 => x"d4",
          8553 => x"d8",
          8554 => x"8c",
          8555 => x"ff",
          8556 => x"82",
          8557 => x"55",
          8558 => x"d8",
          8559 => x"0d",
          8560 => x"0d",
          8561 => x"3d",
          8562 => x"52",
          8563 => x"d7",
          8564 => x"d6",
          8565 => x"82",
          8566 => x"82",
          8567 => x"5e",
          8568 => x"3d",
          8569 => x"cb",
          8570 => x"d6",
          8571 => x"82",
          8572 => x"86",
          8573 => x"82",
          8574 => x"d6",
          8575 => x"2e",
          8576 => x"82",
          8577 => x"80",
          8578 => x"70",
          8579 => x"06",
          8580 => x"54",
          8581 => x"38",
          8582 => x"52",
          8583 => x"52",
          8584 => x"80",
          8585 => x"d8",
          8586 => x"56",
          8587 => x"08",
          8588 => x"54",
          8589 => x"08",
          8590 => x"81",
          8591 => x"82",
          8592 => x"d8",
          8593 => x"09",
          8594 => x"38",
          8595 => x"ba",
          8596 => x"b6",
          8597 => x"d8",
          8598 => x"51",
          8599 => x"3f",
          8600 => x"08",
          8601 => x"d8",
          8602 => x"38",
          8603 => x"52",
          8604 => x"ff",
          8605 => x"78",
          8606 => x"b8",
          8607 => x"54",
          8608 => x"c3",
          8609 => x"88",
          8610 => x"80",
          8611 => x"ff",
          8612 => x"75",
          8613 => x"11",
          8614 => x"b8",
          8615 => x"53",
          8616 => x"53",
          8617 => x"51",
          8618 => x"3f",
          8619 => x"0b",
          8620 => x"34",
          8621 => x"80",
          8622 => x"51",
          8623 => x"3f",
          8624 => x"0b",
          8625 => x"77",
          8626 => x"cd",
          8627 => x"d8",
          8628 => x"d6",
          8629 => x"38",
          8630 => x"0a",
          8631 => x"05",
          8632 => x"ca",
          8633 => x"64",
          8634 => x"ff",
          8635 => x"64",
          8636 => x"8b",
          8637 => x"54",
          8638 => x"15",
          8639 => x"ff",
          8640 => x"82",
          8641 => x"54",
          8642 => x"53",
          8643 => x"51",
          8644 => x"3f",
          8645 => x"d8",
          8646 => x"0d",
          8647 => x"0d",
          8648 => x"05",
          8649 => x"3f",
          8650 => x"3d",
          8651 => x"52",
          8652 => x"d5",
          8653 => x"d6",
          8654 => x"82",
          8655 => x"82",
          8656 => x"4e",
          8657 => x"52",
          8658 => x"52",
          8659 => x"3f",
          8660 => x"08",
          8661 => x"d8",
          8662 => x"38",
          8663 => x"05",
          8664 => x"06",
          8665 => x"73",
          8666 => x"a0",
          8667 => x"08",
          8668 => x"ff",
          8669 => x"ff",
          8670 => x"b0",
          8671 => x"92",
          8672 => x"54",
          8673 => x"3f",
          8674 => x"52",
          8675 => x"d0",
          8676 => x"d8",
          8677 => x"d6",
          8678 => x"38",
          8679 => x"08",
          8680 => x"06",
          8681 => x"a3",
          8682 => x"92",
          8683 => x"81",
          8684 => x"d6",
          8685 => x"2e",
          8686 => x"81",
          8687 => x"51",
          8688 => x"3f",
          8689 => x"08",
          8690 => x"d8",
          8691 => x"38",
          8692 => x"53",
          8693 => x"8d",
          8694 => x"16",
          8695 => x"fd",
          8696 => x"05",
          8697 => x"34",
          8698 => x"70",
          8699 => x"81",
          8700 => x"55",
          8701 => x"74",
          8702 => x"73",
          8703 => x"78",
          8704 => x"83",
          8705 => x"16",
          8706 => x"2a",
          8707 => x"51",
          8708 => x"80",
          8709 => x"38",
          8710 => x"80",
          8711 => x"52",
          8712 => x"b4",
          8713 => x"d6",
          8714 => x"78",
          8715 => x"ee",
          8716 => x"82",
          8717 => x"80",
          8718 => x"38",
          8719 => x"08",
          8720 => x"ff",
          8721 => x"82",
          8722 => x"79",
          8723 => x"58",
          8724 => x"d6",
          8725 => x"c1",
          8726 => x"33",
          8727 => x"2e",
          8728 => x"9a",
          8729 => x"75",
          8730 => x"ff",
          8731 => x"78",
          8732 => x"83",
          8733 => x"39",
          8734 => x"08",
          8735 => x"51",
          8736 => x"82",
          8737 => x"55",
          8738 => x"08",
          8739 => x"51",
          8740 => x"3f",
          8741 => x"08",
          8742 => x"d6",
          8743 => x"3d",
          8744 => x"3d",
          8745 => x"df",
          8746 => x"84",
          8747 => x"05",
          8748 => x"82",
          8749 => x"cc",
          8750 => x"3d",
          8751 => x"3f",
          8752 => x"08",
          8753 => x"d8",
          8754 => x"38",
          8755 => x"52",
          8756 => x"05",
          8757 => x"3f",
          8758 => x"08",
          8759 => x"d8",
          8760 => x"02",
          8761 => x"33",
          8762 => x"54",
          8763 => x"aa",
          8764 => x"06",
          8765 => x"8b",
          8766 => x"06",
          8767 => x"07",
          8768 => x"56",
          8769 => x"34",
          8770 => x"0b",
          8771 => x"78",
          8772 => x"db",
          8773 => x"d8",
          8774 => x"82",
          8775 => x"96",
          8776 => x"ee",
          8777 => x"56",
          8778 => x"3d",
          8779 => x"95",
          8780 => x"92",
          8781 => x"d8",
          8782 => x"d6",
          8783 => x"cb",
          8784 => x"64",
          8785 => x"d0",
          8786 => x"94",
          8787 => x"d8",
          8788 => x"d6",
          8789 => x"38",
          8790 => x"05",
          8791 => x"06",
          8792 => x"73",
          8793 => x"16",
          8794 => x"22",
          8795 => x"07",
          8796 => x"1f",
          8797 => x"b6",
          8798 => x"81",
          8799 => x"34",
          8800 => x"a1",
          8801 => x"d6",
          8802 => x"74",
          8803 => x"0c",
          8804 => x"04",
          8805 => x"6a",
          8806 => x"80",
          8807 => x"cc",
          8808 => x"3d",
          8809 => x"3f",
          8810 => x"08",
          8811 => x"08",
          8812 => x"d6",
          8813 => x"80",
          8814 => x"57",
          8815 => x"81",
          8816 => x"70",
          8817 => x"55",
          8818 => x"80",
          8819 => x"5d",
          8820 => x"52",
          8821 => x"52",
          8822 => x"db",
          8823 => x"d8",
          8824 => x"d6",
          8825 => x"d2",
          8826 => x"73",
          8827 => x"bc",
          8828 => x"d8",
          8829 => x"d6",
          8830 => x"38",
          8831 => x"08",
          8832 => x"08",
          8833 => x"56",
          8834 => x"19",
          8835 => x"59",
          8836 => x"74",
          8837 => x"56",
          8838 => x"ec",
          8839 => x"75",
          8840 => x"74",
          8841 => x"2e",
          8842 => x"16",
          8843 => x"33",
          8844 => x"73",
          8845 => x"38",
          8846 => x"84",
          8847 => x"06",
          8848 => x"7a",
          8849 => x"76",
          8850 => x"07",
          8851 => x"54",
          8852 => x"80",
          8853 => x"80",
          8854 => x"7b",
          8855 => x"53",
          8856 => x"c4",
          8857 => x"d8",
          8858 => x"d6",
          8859 => x"38",
          8860 => x"55",
          8861 => x"56",
          8862 => x"8b",
          8863 => x"56",
          8864 => x"83",
          8865 => x"75",
          8866 => x"51",
          8867 => x"3f",
          8868 => x"08",
          8869 => x"82",
          8870 => x"99",
          8871 => x"e6",
          8872 => x"53",
          8873 => x"b4",
          8874 => x"3d",
          8875 => x"3f",
          8876 => x"08",
          8877 => x"08",
          8878 => x"d6",
          8879 => x"dd",
          8880 => x"a0",
          8881 => x"70",
          8882 => x"9c",
          8883 => x"6d",
          8884 => x"55",
          8885 => x"27",
          8886 => x"77",
          8887 => x"51",
          8888 => x"3f",
          8889 => x"08",
          8890 => x"26",
          8891 => x"82",
          8892 => x"51",
          8893 => x"83",
          8894 => x"d6",
          8895 => x"93",
          8896 => x"d6",
          8897 => x"ff",
          8898 => x"74",
          8899 => x"38",
          8900 => x"c8",
          8901 => x"9c",
          8902 => x"d6",
          8903 => x"38",
          8904 => x"27",
          8905 => x"89",
          8906 => x"8b",
          8907 => x"27",
          8908 => x"55",
          8909 => x"81",
          8910 => x"8f",
          8911 => x"2a",
          8912 => x"70",
          8913 => x"34",
          8914 => x"74",
          8915 => x"05",
          8916 => x"16",
          8917 => x"51",
          8918 => x"9f",
          8919 => x"38",
          8920 => x"54",
          8921 => x"81",
          8922 => x"b1",
          8923 => x"2e",
          8924 => x"a3",
          8925 => x"15",
          8926 => x"54",
          8927 => x"09",
          8928 => x"38",
          8929 => x"75",
          8930 => x"40",
          8931 => x"52",
          8932 => x"52",
          8933 => x"9f",
          8934 => x"d8",
          8935 => x"d6",
          8936 => x"f7",
          8937 => x"74",
          8938 => x"80",
          8939 => x"d8",
          8940 => x"d6",
          8941 => x"38",
          8942 => x"38",
          8943 => x"74",
          8944 => x"39",
          8945 => x"08",
          8946 => x"81",
          8947 => x"38",
          8948 => x"74",
          8949 => x"38",
          8950 => x"51",
          8951 => x"3f",
          8952 => x"08",
          8953 => x"d8",
          8954 => x"a0",
          8955 => x"d8",
          8956 => x"51",
          8957 => x"3f",
          8958 => x"0b",
          8959 => x"8b",
          8960 => x"66",
          8961 => x"d5",
          8962 => x"81",
          8963 => x"34",
          8964 => x"9c",
          8965 => x"d6",
          8966 => x"73",
          8967 => x"d6",
          8968 => x"3d",
          8969 => x"3d",
          8970 => x"02",
          8971 => x"cb",
          8972 => x"3d",
          8973 => x"72",
          8974 => x"5a",
          8975 => x"82",
          8976 => x"58",
          8977 => x"08",
          8978 => x"91",
          8979 => x"77",
          8980 => x"7c",
          8981 => x"38",
          8982 => x"59",
          8983 => x"90",
          8984 => x"81",
          8985 => x"06",
          8986 => x"73",
          8987 => x"54",
          8988 => x"82",
          8989 => x"39",
          8990 => x"8b",
          8991 => x"11",
          8992 => x"2b",
          8993 => x"54",
          8994 => x"fe",
          8995 => x"ff",
          8996 => x"70",
          8997 => x"07",
          8998 => x"d6",
          8999 => x"90",
          9000 => x"40",
          9001 => x"55",
          9002 => x"88",
          9003 => x"08",
          9004 => x"38",
          9005 => x"77",
          9006 => x"56",
          9007 => x"51",
          9008 => x"3f",
          9009 => x"55",
          9010 => x"08",
          9011 => x"38",
          9012 => x"d6",
          9013 => x"2e",
          9014 => x"82",
          9015 => x"ff",
          9016 => x"38",
          9017 => x"08",
          9018 => x"16",
          9019 => x"2e",
          9020 => x"87",
          9021 => x"74",
          9022 => x"74",
          9023 => x"81",
          9024 => x"38",
          9025 => x"ff",
          9026 => x"2e",
          9027 => x"7b",
          9028 => x"80",
          9029 => x"81",
          9030 => x"81",
          9031 => x"06",
          9032 => x"56",
          9033 => x"52",
          9034 => x"9e",
          9035 => x"d6",
          9036 => x"82",
          9037 => x"80",
          9038 => x"81",
          9039 => x"56",
          9040 => x"d3",
          9041 => x"ff",
          9042 => x"7c",
          9043 => x"55",
          9044 => x"b3",
          9045 => x"1b",
          9046 => x"1b",
          9047 => x"33",
          9048 => x"54",
          9049 => x"34",
          9050 => x"fe",
          9051 => x"08",
          9052 => x"74",
          9053 => x"75",
          9054 => x"16",
          9055 => x"33",
          9056 => x"73",
          9057 => x"77",
          9058 => x"d6",
          9059 => x"3d",
          9060 => x"3d",
          9061 => x"02",
          9062 => x"eb",
          9063 => x"3d",
          9064 => x"59",
          9065 => x"8b",
          9066 => x"82",
          9067 => x"24",
          9068 => x"82",
          9069 => x"84",
          9070 => x"a0",
          9071 => x"51",
          9072 => x"2e",
          9073 => x"75",
          9074 => x"d8",
          9075 => x"06",
          9076 => x"7e",
          9077 => x"fe",
          9078 => x"d8",
          9079 => x"06",
          9080 => x"56",
          9081 => x"74",
          9082 => x"76",
          9083 => x"81",
          9084 => x"8a",
          9085 => x"b2",
          9086 => x"fc",
          9087 => x"52",
          9088 => x"93",
          9089 => x"d6",
          9090 => x"38",
          9091 => x"80",
          9092 => x"74",
          9093 => x"26",
          9094 => x"15",
          9095 => x"74",
          9096 => x"38",
          9097 => x"80",
          9098 => x"84",
          9099 => x"92",
          9100 => x"80",
          9101 => x"38",
          9102 => x"06",
          9103 => x"2e",
          9104 => x"56",
          9105 => x"78",
          9106 => x"89",
          9107 => x"2b",
          9108 => x"43",
          9109 => x"38",
          9110 => x"30",
          9111 => x"77",
          9112 => x"91",
          9113 => x"c2",
          9114 => x"f8",
          9115 => x"52",
          9116 => x"92",
          9117 => x"56",
          9118 => x"08",
          9119 => x"77",
          9120 => x"77",
          9121 => x"d8",
          9122 => x"45",
          9123 => x"bf",
          9124 => x"8e",
          9125 => x"26",
          9126 => x"74",
          9127 => x"48",
          9128 => x"75",
          9129 => x"38",
          9130 => x"81",
          9131 => x"fa",
          9132 => x"2a",
          9133 => x"56",
          9134 => x"2e",
          9135 => x"87",
          9136 => x"82",
          9137 => x"38",
          9138 => x"55",
          9139 => x"83",
          9140 => x"81",
          9141 => x"56",
          9142 => x"80",
          9143 => x"38",
          9144 => x"83",
          9145 => x"06",
          9146 => x"78",
          9147 => x"91",
          9148 => x"0b",
          9149 => x"22",
          9150 => x"80",
          9151 => x"74",
          9152 => x"38",
          9153 => x"56",
          9154 => x"17",
          9155 => x"57",
          9156 => x"2e",
          9157 => x"75",
          9158 => x"79",
          9159 => x"fe",
          9160 => x"82",
          9161 => x"84",
          9162 => x"05",
          9163 => x"5e",
          9164 => x"80",
          9165 => x"d8",
          9166 => x"8a",
          9167 => x"fd",
          9168 => x"75",
          9169 => x"38",
          9170 => x"78",
          9171 => x"8c",
          9172 => x"0b",
          9173 => x"22",
          9174 => x"80",
          9175 => x"74",
          9176 => x"38",
          9177 => x"56",
          9178 => x"17",
          9179 => x"57",
          9180 => x"2e",
          9181 => x"75",
          9182 => x"79",
          9183 => x"fe",
          9184 => x"82",
          9185 => x"10",
          9186 => x"82",
          9187 => x"9f",
          9188 => x"38",
          9189 => x"d6",
          9190 => x"82",
          9191 => x"05",
          9192 => x"2a",
          9193 => x"56",
          9194 => x"17",
          9195 => x"81",
          9196 => x"60",
          9197 => x"65",
          9198 => x"12",
          9199 => x"30",
          9200 => x"74",
          9201 => x"59",
          9202 => x"7d",
          9203 => x"81",
          9204 => x"76",
          9205 => x"41",
          9206 => x"76",
          9207 => x"90",
          9208 => x"62",
          9209 => x"51",
          9210 => x"26",
          9211 => x"75",
          9212 => x"31",
          9213 => x"65",
          9214 => x"fe",
          9215 => x"82",
          9216 => x"58",
          9217 => x"09",
          9218 => x"38",
          9219 => x"08",
          9220 => x"26",
          9221 => x"78",
          9222 => x"79",
          9223 => x"78",
          9224 => x"86",
          9225 => x"82",
          9226 => x"06",
          9227 => x"83",
          9228 => x"82",
          9229 => x"27",
          9230 => x"8f",
          9231 => x"55",
          9232 => x"26",
          9233 => x"59",
          9234 => x"62",
          9235 => x"74",
          9236 => x"38",
          9237 => x"88",
          9238 => x"d8",
          9239 => x"26",
          9240 => x"86",
          9241 => x"1a",
          9242 => x"79",
          9243 => x"38",
          9244 => x"80",
          9245 => x"2e",
          9246 => x"83",
          9247 => x"9f",
          9248 => x"8b",
          9249 => x"06",
          9250 => x"74",
          9251 => x"84",
          9252 => x"52",
          9253 => x"90",
          9254 => x"53",
          9255 => x"52",
          9256 => x"90",
          9257 => x"80",
          9258 => x"51",
          9259 => x"3f",
          9260 => x"34",
          9261 => x"ff",
          9262 => x"1b",
          9263 => x"d0",
          9264 => x"90",
          9265 => x"83",
          9266 => x"70",
          9267 => x"80",
          9268 => x"55",
          9269 => x"ff",
          9270 => x"66",
          9271 => x"ff",
          9272 => x"38",
          9273 => x"ff",
          9274 => x"1b",
          9275 => x"a0",
          9276 => x"74",
          9277 => x"51",
          9278 => x"3f",
          9279 => x"1c",
          9280 => x"98",
          9281 => x"8f",
          9282 => x"ff",
          9283 => x"51",
          9284 => x"3f",
          9285 => x"1b",
          9286 => x"92",
          9287 => x"2e",
          9288 => x"80",
          9289 => x"88",
          9290 => x"80",
          9291 => x"ff",
          9292 => x"7c",
          9293 => x"51",
          9294 => x"3f",
          9295 => x"1b",
          9296 => x"ea",
          9297 => x"b0",
          9298 => x"8e",
          9299 => x"52",
          9300 => x"ff",
          9301 => x"ff",
          9302 => x"c0",
          9303 => x"0b",
          9304 => x"34",
          9305 => x"c7",
          9306 => x"c7",
          9307 => x"39",
          9308 => x"0a",
          9309 => x"51",
          9310 => x"3f",
          9311 => x"ff",
          9312 => x"1b",
          9313 => x"88",
          9314 => x"0b",
          9315 => x"a9",
          9316 => x"34",
          9317 => x"c7",
          9318 => x"1b",
          9319 => x"bd",
          9320 => x"d5",
          9321 => x"1b",
          9322 => x"ff",
          9323 => x"81",
          9324 => x"7a",
          9325 => x"ff",
          9326 => x"81",
          9327 => x"d8",
          9328 => x"38",
          9329 => x"09",
          9330 => x"ee",
          9331 => x"60",
          9332 => x"7a",
          9333 => x"ff",
          9334 => x"84",
          9335 => x"52",
          9336 => x"8e",
          9337 => x"8b",
          9338 => x"52",
          9339 => x"8d",
          9340 => x"8a",
          9341 => x"52",
          9342 => x"51",
          9343 => x"3f",
          9344 => x"83",
          9345 => x"ff",
          9346 => x"82",
          9347 => x"1b",
          9348 => x"9a",
          9349 => x"d5",
          9350 => x"ff",
          9351 => x"75",
          9352 => x"05",
          9353 => x"7e",
          9354 => x"93",
          9355 => x"60",
          9356 => x"52",
          9357 => x"89",
          9358 => x"53",
          9359 => x"51",
          9360 => x"3f",
          9361 => x"58",
          9362 => x"09",
          9363 => x"38",
          9364 => x"51",
          9365 => x"3f",
          9366 => x"1b",
          9367 => x"ce",
          9368 => x"52",
          9369 => x"91",
          9370 => x"ff",
          9371 => x"81",
          9372 => x"f8",
          9373 => x"7a",
          9374 => x"b2",
          9375 => x"61",
          9376 => x"26",
          9377 => x"57",
          9378 => x"53",
          9379 => x"51",
          9380 => x"3f",
          9381 => x"08",
          9382 => x"84",
          9383 => x"d6",
          9384 => x"7a",
          9385 => x"d8",
          9386 => x"75",
          9387 => x"56",
          9388 => x"81",
          9389 => x"80",
          9390 => x"38",
          9391 => x"83",
          9392 => x"63",
          9393 => x"74",
          9394 => x"38",
          9395 => x"54",
          9396 => x"52",
          9397 => x"87",
          9398 => x"d6",
          9399 => x"c1",
          9400 => x"75",
          9401 => x"56",
          9402 => x"8c",
          9403 => x"2e",
          9404 => x"56",
          9405 => x"ff",
          9406 => x"84",
          9407 => x"2e",
          9408 => x"56",
          9409 => x"58",
          9410 => x"38",
          9411 => x"77",
          9412 => x"ff",
          9413 => x"82",
          9414 => x"78",
          9415 => x"f0",
          9416 => x"1b",
          9417 => x"34",
          9418 => x"16",
          9419 => x"82",
          9420 => x"83",
          9421 => x"84",
          9422 => x"67",
          9423 => x"fd",
          9424 => x"51",
          9425 => x"3f",
          9426 => x"16",
          9427 => x"d8",
          9428 => x"bf",
          9429 => x"86",
          9430 => x"d6",
          9431 => x"16",
          9432 => x"83",
          9433 => x"ff",
          9434 => x"66",
          9435 => x"1b",
          9436 => x"ba",
          9437 => x"77",
          9438 => x"7e",
          9439 => x"bf",
          9440 => x"82",
          9441 => x"a2",
          9442 => x"80",
          9443 => x"ff",
          9444 => x"81",
          9445 => x"d8",
          9446 => x"89",
          9447 => x"8a",
          9448 => x"86",
          9449 => x"d8",
          9450 => x"82",
          9451 => x"99",
          9452 => x"f5",
          9453 => x"60",
          9454 => x"79",
          9455 => x"5a",
          9456 => x"78",
          9457 => x"8d",
          9458 => x"55",
          9459 => x"fc",
          9460 => x"51",
          9461 => x"7a",
          9462 => x"81",
          9463 => x"8c",
          9464 => x"74",
          9465 => x"38",
          9466 => x"81",
          9467 => x"81",
          9468 => x"8a",
          9469 => x"06",
          9470 => x"76",
          9471 => x"76",
          9472 => x"55",
          9473 => x"d8",
          9474 => x"0d",
          9475 => x"0d",
          9476 => x"05",
          9477 => x"59",
          9478 => x"2e",
          9479 => x"87",
          9480 => x"76",
          9481 => x"84",
          9482 => x"80",
          9483 => x"38",
          9484 => x"77",
          9485 => x"56",
          9486 => x"34",
          9487 => x"bb",
          9488 => x"38",
          9489 => x"05",
          9490 => x"8c",
          9491 => x"08",
          9492 => x"3f",
          9493 => x"70",
          9494 => x"07",
          9495 => x"30",
          9496 => x"56",
          9497 => x"0c",
          9498 => x"18",
          9499 => x"0d",
          9500 => x"0d",
          9501 => x"08",
          9502 => x"75",
          9503 => x"89",
          9504 => x"54",
          9505 => x"16",
          9506 => x"51",
          9507 => x"82",
          9508 => x"91",
          9509 => x"08",
          9510 => x"81",
          9511 => x"88",
          9512 => x"83",
          9513 => x"74",
          9514 => x"0c",
          9515 => x"04",
          9516 => x"75",
          9517 => x"53",
          9518 => x"51",
          9519 => x"3f",
          9520 => x"85",
          9521 => x"ea",
          9522 => x"80",
          9523 => x"6a",
          9524 => x"70",
          9525 => x"d8",
          9526 => x"72",
          9527 => x"3f",
          9528 => x"8d",
          9529 => x"0d",
          9530 => x"0d",
          9531 => x"05",
          9532 => x"55",
          9533 => x"72",
          9534 => x"8a",
          9535 => x"ff",
          9536 => x"80",
          9537 => x"ff",
          9538 => x"51",
          9539 => x"2e",
          9540 => x"b4",
          9541 => x"2e",
          9542 => x"c9",
          9543 => x"72",
          9544 => x"38",
          9545 => x"83",
          9546 => x"53",
          9547 => x"ff",
          9548 => x"71",
          9549 => x"98",
          9550 => x"51",
          9551 => x"81",
          9552 => x"81",
          9553 => x"51",
          9554 => x"d8",
          9555 => x"0d",
          9556 => x"0d",
          9557 => x"22",
          9558 => x"96",
          9559 => x"51",
          9560 => x"80",
          9561 => x"38",
          9562 => x"39",
          9563 => x"2e",
          9564 => x"91",
          9565 => x"ff",
          9566 => x"70",
          9567 => x"98",
          9568 => x"54",
          9569 => x"d6",
          9570 => x"3d",
          9571 => x"3d",
          9572 => x"70",
          9573 => x"26",
          9574 => x"70",
          9575 => x"06",
          9576 => x"57",
          9577 => x"72",
          9578 => x"82",
          9579 => x"75",
          9580 => x"57",
          9581 => x"70",
          9582 => x"75",
          9583 => x"52",
          9584 => x"fb",
          9585 => x"82",
          9586 => x"70",
          9587 => x"81",
          9588 => x"18",
          9589 => x"53",
          9590 => x"80",
          9591 => x"88",
          9592 => x"38",
          9593 => x"82",
          9594 => x"51",
          9595 => x"71",
          9596 => x"76",
          9597 => x"54",
          9598 => x"c3",
          9599 => x"31",
          9600 => x"71",
          9601 => x"a4",
          9602 => x"51",
          9603 => x"12",
          9604 => x"d0",
          9605 => x"39",
          9606 => x"90",
          9607 => x"51",
          9608 => x"b0",
          9609 => x"39",
          9610 => x"51",
          9611 => x"ff",
          9612 => x"39",
          9613 => x"38",
          9614 => x"56",
          9615 => x"71",
          9616 => x"d6",
          9617 => x"3d",
          9618 => x"00",
          9619 => x"ff",
          9620 => x"ff",
          9621 => x"00",
          9622 => x"ff",
          9623 => x"2c",
          9624 => x"2b",
          9625 => x"2b",
          9626 => x"2b",
          9627 => x"2b",
          9628 => x"2b",
          9629 => x"2b",
          9630 => x"2b",
          9631 => x"2c",
          9632 => x"2c",
          9633 => x"2c",
          9634 => x"2c",
          9635 => x"2c",
          9636 => x"2c",
          9637 => x"2c",
          9638 => x"2c",
          9639 => x"2c",
          9640 => x"2c",
          9641 => x"2c",
          9642 => x"2c",
          9643 => x"42",
          9644 => x"42",
          9645 => x"42",
          9646 => x"42",
          9647 => x"42",
          9648 => x"48",
          9649 => x"49",
          9650 => x"4a",
          9651 => x"4c",
          9652 => x"49",
          9653 => x"46",
          9654 => x"4b",
          9655 => x"4c",
          9656 => x"4b",
          9657 => x"4b",
          9658 => x"4b",
          9659 => x"49",
          9660 => x"46",
          9661 => x"4a",
          9662 => x"4a",
          9663 => x"4b",
          9664 => x"46",
          9665 => x"46",
          9666 => x"4b",
          9667 => x"4b",
          9668 => x"4c",
          9669 => x"4c",
          9670 => x"95",
          9671 => x"95",
          9672 => x"96",
          9673 => x"96",
          9674 => x"96",
          9675 => x"96",
          9676 => x"96",
          9677 => x"96",
          9678 => x"96",
          9679 => x"0e",
          9680 => x"17",
          9681 => x"17",
          9682 => x"0e",
          9683 => x"17",
          9684 => x"17",
          9685 => x"17",
          9686 => x"17",
          9687 => x"17",
          9688 => x"17",
          9689 => x"17",
          9690 => x"0e",
          9691 => x"17",
          9692 => x"0e",
          9693 => x"0e",
          9694 => x"17",
          9695 => x"17",
          9696 => x"17",
          9697 => x"17",
          9698 => x"17",
          9699 => x"17",
          9700 => x"17",
          9701 => x"17",
          9702 => x"17",
          9703 => x"17",
          9704 => x"17",
          9705 => x"17",
          9706 => x"17",
          9707 => x"17",
          9708 => x"17",
          9709 => x"17",
          9710 => x"17",
          9711 => x"17",
          9712 => x"17",
          9713 => x"17",
          9714 => x"17",
          9715 => x"17",
          9716 => x"17",
          9717 => x"17",
          9718 => x"17",
          9719 => x"17",
          9720 => x"17",
          9721 => x"17",
          9722 => x"17",
          9723 => x"17",
          9724 => x"17",
          9725 => x"17",
          9726 => x"17",
          9727 => x"17",
          9728 => x"17",
          9729 => x"17",
          9730 => x"0f",
          9731 => x"17",
          9732 => x"17",
          9733 => x"17",
          9734 => x"17",
          9735 => x"11",
          9736 => x"17",
          9737 => x"17",
          9738 => x"17",
          9739 => x"17",
          9740 => x"17",
          9741 => x"17",
          9742 => x"17",
          9743 => x"17",
          9744 => x"17",
          9745 => x"17",
          9746 => x"0e",
          9747 => x"10",
          9748 => x"0e",
          9749 => x"0e",
          9750 => x"0e",
          9751 => x"17",
          9752 => x"10",
          9753 => x"17",
          9754 => x"17",
          9755 => x"0e",
          9756 => x"17",
          9757 => x"17",
          9758 => x"10",
          9759 => x"10",
          9760 => x"17",
          9761 => x"17",
          9762 => x"0f",
          9763 => x"17",
          9764 => x"11",
          9765 => x"17",
          9766 => x"17",
          9767 => x"11",
          9768 => x"6e",
          9769 => x"00",
          9770 => x"6f",
          9771 => x"00",
          9772 => x"6e",
          9773 => x"00",
          9774 => x"6f",
          9775 => x"00",
          9776 => x"78",
          9777 => x"00",
          9778 => x"6c",
          9779 => x"00",
          9780 => x"6f",
          9781 => x"00",
          9782 => x"69",
          9783 => x"00",
          9784 => x"75",
          9785 => x"00",
          9786 => x"62",
          9787 => x"68",
          9788 => x"77",
          9789 => x"64",
          9790 => x"65",
          9791 => x"64",
          9792 => x"65",
          9793 => x"6c",
          9794 => x"00",
          9795 => x"70",
          9796 => x"73",
          9797 => x"74",
          9798 => x"73",
          9799 => x"00",
          9800 => x"66",
          9801 => x"00",
          9802 => x"73",
          9803 => x"00",
          9804 => x"61",
          9805 => x"00",
          9806 => x"61",
          9807 => x"00",
          9808 => x"6c",
          9809 => x"00",
          9810 => x"00",
          9811 => x"73",
          9812 => x"72",
          9813 => x"00",
          9814 => x"74",
          9815 => x"61",
          9816 => x"72",
          9817 => x"2e",
          9818 => x"73",
          9819 => x"6f",
          9820 => x"65",
          9821 => x"2e",
          9822 => x"20",
          9823 => x"65",
          9824 => x"75",
          9825 => x"00",
          9826 => x"20",
          9827 => x"68",
          9828 => x"75",
          9829 => x"00",
          9830 => x"76",
          9831 => x"64",
          9832 => x"6c",
          9833 => x"6d",
          9834 => x"00",
          9835 => x"63",
          9836 => x"20",
          9837 => x"69",
          9838 => x"00",
          9839 => x"6c",
          9840 => x"6c",
          9841 => x"64",
          9842 => x"78",
          9843 => x"73",
          9844 => x"00",
          9845 => x"6c",
          9846 => x"61",
          9847 => x"65",
          9848 => x"76",
          9849 => x"64",
          9850 => x"00",
          9851 => x"20",
          9852 => x"77",
          9853 => x"65",
          9854 => x"6f",
          9855 => x"74",
          9856 => x"00",
          9857 => x"69",
          9858 => x"6e",
          9859 => x"65",
          9860 => x"73",
          9861 => x"76",
          9862 => x"64",
          9863 => x"00",
          9864 => x"73",
          9865 => x"6f",
          9866 => x"6e",
          9867 => x"65",
          9868 => x"00",
          9869 => x"20",
          9870 => x"70",
          9871 => x"62",
          9872 => x"66",
          9873 => x"73",
          9874 => x"65",
          9875 => x"6f",
          9876 => x"20",
          9877 => x"64",
          9878 => x"2e",
          9879 => x"72",
          9880 => x"20",
          9881 => x"72",
          9882 => x"2e",
          9883 => x"6d",
          9884 => x"74",
          9885 => x"70",
          9886 => x"74",
          9887 => x"20",
          9888 => x"63",
          9889 => x"65",
          9890 => x"00",
          9891 => x"6c",
          9892 => x"73",
          9893 => x"63",
          9894 => x"2e",
          9895 => x"73",
          9896 => x"69",
          9897 => x"6e",
          9898 => x"65",
          9899 => x"79",
          9900 => x"00",
          9901 => x"6f",
          9902 => x"6e",
          9903 => x"70",
          9904 => x"66",
          9905 => x"73",
          9906 => x"00",
          9907 => x"72",
          9908 => x"74",
          9909 => x"20",
          9910 => x"6f",
          9911 => x"63",
          9912 => x"00",
          9913 => x"63",
          9914 => x"73",
          9915 => x"00",
          9916 => x"6b",
          9917 => x"6e",
          9918 => x"72",
          9919 => x"00",
          9920 => x"6c",
          9921 => x"79",
          9922 => x"20",
          9923 => x"61",
          9924 => x"6c",
          9925 => x"79",
          9926 => x"2f",
          9927 => x"2e",
          9928 => x"00",
          9929 => x"61",
          9930 => x"00",
          9931 => x"25",
          9932 => x"78",
          9933 => x"3d",
          9934 => x"6c",
          9935 => x"32",
          9936 => x"38",
          9937 => x"20",
          9938 => x"42",
          9939 => x"38",
          9940 => x"25",
          9941 => x"78",
          9942 => x"38",
          9943 => x"00",
          9944 => x"38",
          9945 => x"00",
          9946 => x"20",
          9947 => x"34",
          9948 => x"00",
          9949 => x"20",
          9950 => x"20",
          9951 => x"00",
          9952 => x"32",
          9953 => x"00",
          9954 => x"00",
          9955 => x"00",
          9956 => x"00",
          9957 => x"53",
          9958 => x"2a",
          9959 => x"20",
          9960 => x"00",
          9961 => x"2f",
          9962 => x"32",
          9963 => x"00",
          9964 => x"2e",
          9965 => x"00",
          9966 => x"50",
          9967 => x"72",
          9968 => x"25",
          9969 => x"29",
          9970 => x"20",
          9971 => x"2a",
          9972 => x"00",
          9973 => x"55",
          9974 => x"74",
          9975 => x"75",
          9976 => x"48",
          9977 => x"6c",
          9978 => x"00",
          9979 => x"6d",
          9980 => x"69",
          9981 => x"72",
          9982 => x"74",
          9983 => x"32",
          9984 => x"74",
          9985 => x"75",
          9986 => x"00",
          9987 => x"43",
          9988 => x"52",
          9989 => x"6e",
          9990 => x"72",
          9991 => x"00",
          9992 => x"43",
          9993 => x"57",
          9994 => x"6e",
          9995 => x"72",
          9996 => x"00",
          9997 => x"52",
          9998 => x"52",
          9999 => x"6e",
         10000 => x"72",
         10001 => x"00",
         10002 => x"52",
         10003 => x"54",
         10004 => x"6e",
         10005 => x"72",
         10006 => x"00",
         10007 => x"52",
         10008 => x"52",
         10009 => x"6e",
         10010 => x"72",
         10011 => x"00",
         10012 => x"52",
         10013 => x"54",
         10014 => x"6e",
         10015 => x"72",
         10016 => x"00",
         10017 => x"74",
         10018 => x"67",
         10019 => x"20",
         10020 => x"65",
         10021 => x"2e",
         10022 => x"61",
         10023 => x"6e",
         10024 => x"69",
         10025 => x"2e",
         10026 => x"00",
         10027 => x"74",
         10028 => x"65",
         10029 => x"61",
         10030 => x"00",
         10031 => x"53",
         10032 => x"74",
         10033 => x"00",
         10034 => x"69",
         10035 => x"20",
         10036 => x"69",
         10037 => x"69",
         10038 => x"73",
         10039 => x"64",
         10040 => x"72",
         10041 => x"2c",
         10042 => x"65",
         10043 => x"20",
         10044 => x"74",
         10045 => x"6e",
         10046 => x"6c",
         10047 => x"00",
         10048 => x"00",
         10049 => x"65",
         10050 => x"6e",
         10051 => x"2e",
         10052 => x"00",
         10053 => x"70",
         10054 => x"67",
         10055 => x"00",
         10056 => x"6d",
         10057 => x"69",
         10058 => x"2e",
         10059 => x"00",
         10060 => x"38",
         10061 => x"25",
         10062 => x"29",
         10063 => x"30",
         10064 => x"28",
         10065 => x"78",
         10066 => x"00",
         10067 => x"6d",
         10068 => x"65",
         10069 => x"79",
         10070 => x"6f",
         10071 => x"65",
         10072 => x"00",
         10073 => x"38",
         10074 => x"25",
         10075 => x"2d",
         10076 => x"3f",
         10077 => x"38",
         10078 => x"25",
         10079 => x"2d",
         10080 => x"38",
         10081 => x"25",
         10082 => x"58",
         10083 => x"00",
         10084 => x"65",
         10085 => x"69",
         10086 => x"63",
         10087 => x"20",
         10088 => x"30",
         10089 => x"20",
         10090 => x"0a",
         10091 => x"6c",
         10092 => x"67",
         10093 => x"64",
         10094 => x"20",
         10095 => x"6c",
         10096 => x"2e",
         10097 => x"00",
         10098 => x"6c",
         10099 => x"65",
         10100 => x"6e",
         10101 => x"63",
         10102 => x"20",
         10103 => x"29",
         10104 => x"00",
         10105 => x"73",
         10106 => x"74",
         10107 => x"20",
         10108 => x"6c",
         10109 => x"74",
         10110 => x"2e",
         10111 => x"00",
         10112 => x"6c",
         10113 => x"65",
         10114 => x"74",
         10115 => x"2e",
         10116 => x"00",
         10117 => x"55",
         10118 => x"6e",
         10119 => x"3a",
         10120 => x"5c",
         10121 => x"25",
         10122 => x"00",
         10123 => x"3a",
         10124 => x"5c",
         10125 => x"00",
         10126 => x"3a",
         10127 => x"00",
         10128 => x"64",
         10129 => x"6d",
         10130 => x"64",
         10131 => x"00",
         10132 => x"6d",
         10133 => x"20",
         10134 => x"61",
         10135 => x"65",
         10136 => x"63",
         10137 => x"6f",
         10138 => x"72",
         10139 => x"73",
         10140 => x"6f",
         10141 => x"6e",
         10142 => x"00",
         10143 => x"73",
         10144 => x"67",
         10145 => x"69",
         10146 => x"00",
         10147 => x"6e",
         10148 => x"67",
         10149 => x"00",
         10150 => x"61",
         10151 => x"6e",
         10152 => x"6e",
         10153 => x"72",
         10154 => x"73",
         10155 => x"00",
         10156 => x"2f",
         10157 => x"25",
         10158 => x"64",
         10159 => x"3a",
         10160 => x"25",
         10161 => x"0a",
         10162 => x"43",
         10163 => x"6e",
         10164 => x"75",
         10165 => x"69",
         10166 => x"00",
         10167 => x"66",
         10168 => x"20",
         10169 => x"20",
         10170 => x"66",
         10171 => x"00",
         10172 => x"44",
         10173 => x"63",
         10174 => x"69",
         10175 => x"65",
         10176 => x"74",
         10177 => x"00",
         10178 => x"20",
         10179 => x"20",
         10180 => x"41",
         10181 => x"28",
         10182 => x"58",
         10183 => x"38",
         10184 => x"0a",
         10185 => x"20",
         10186 => x"52",
         10187 => x"20",
         10188 => x"28",
         10189 => x"58",
         10190 => x"38",
         10191 => x"0a",
         10192 => x"20",
         10193 => x"53",
         10194 => x"52",
         10195 => x"28",
         10196 => x"58",
         10197 => x"38",
         10198 => x"0a",
         10199 => x"20",
         10200 => x"41",
         10201 => x"20",
         10202 => x"28",
         10203 => x"58",
         10204 => x"38",
         10205 => x"0a",
         10206 => x"20",
         10207 => x"4d",
         10208 => x"20",
         10209 => x"28",
         10210 => x"58",
         10211 => x"38",
         10212 => x"0a",
         10213 => x"20",
         10214 => x"20",
         10215 => x"44",
         10216 => x"28",
         10217 => x"69",
         10218 => x"20",
         10219 => x"32",
         10220 => x"0a",
         10221 => x"20",
         10222 => x"4d",
         10223 => x"20",
         10224 => x"28",
         10225 => x"65",
         10226 => x"20",
         10227 => x"32",
         10228 => x"0a",
         10229 => x"20",
         10230 => x"54",
         10231 => x"54",
         10232 => x"28",
         10233 => x"6e",
         10234 => x"73",
         10235 => x"32",
         10236 => x"0a",
         10237 => x"20",
         10238 => x"53",
         10239 => x"4e",
         10240 => x"55",
         10241 => x"00",
         10242 => x"20",
         10243 => x"20",
         10244 => x"00",
         10245 => x"20",
         10246 => x"43",
         10247 => x"00",
         10248 => x"20",
         10249 => x"32",
         10250 => x"20",
         10251 => x"49",
         10252 => x"64",
         10253 => x"73",
         10254 => x"00",
         10255 => x"20",
         10256 => x"55",
         10257 => x"73",
         10258 => x"56",
         10259 => x"6f",
         10260 => x"64",
         10261 => x"73",
         10262 => x"20",
         10263 => x"58",
         10264 => x"00",
         10265 => x"20",
         10266 => x"55",
         10267 => x"6d",
         10268 => x"20",
         10269 => x"72",
         10270 => x"64",
         10271 => x"73",
         10272 => x"20",
         10273 => x"58",
         10274 => x"00",
         10275 => x"20",
         10276 => x"61",
         10277 => x"53",
         10278 => x"74",
         10279 => x"64",
         10280 => x"73",
         10281 => x"20",
         10282 => x"20",
         10283 => x"58",
         10284 => x"00",
         10285 => x"73",
         10286 => x"00",
         10287 => x"20",
         10288 => x"55",
         10289 => x"20",
         10290 => x"20",
         10291 => x"20",
         10292 => x"20",
         10293 => x"20",
         10294 => x"20",
         10295 => x"58",
         10296 => x"00",
         10297 => x"20",
         10298 => x"73",
         10299 => x"20",
         10300 => x"63",
         10301 => x"72",
         10302 => x"20",
         10303 => x"20",
         10304 => x"20",
         10305 => x"25",
         10306 => x"4d",
         10307 => x"00",
         10308 => x"20",
         10309 => x"52",
         10310 => x"43",
         10311 => x"6b",
         10312 => x"65",
         10313 => x"20",
         10314 => x"20",
         10315 => x"20",
         10316 => x"25",
         10317 => x"4d",
         10318 => x"00",
         10319 => x"20",
         10320 => x"73",
         10321 => x"6e",
         10322 => x"44",
         10323 => x"20",
         10324 => x"63",
         10325 => x"72",
         10326 => x"20",
         10327 => x"25",
         10328 => x"4d",
         10329 => x"00",
         10330 => x"61",
         10331 => x"00",
         10332 => x"64",
         10333 => x"00",
         10334 => x"65",
         10335 => x"00",
         10336 => x"4f",
         10337 => x"4f",
         10338 => x"00",
         10339 => x"6b",
         10340 => x"6e",
         10341 => x"a2",
         10342 => x"00",
         10343 => x"00",
         10344 => x"a2",
         10345 => x"00",
         10346 => x"00",
         10347 => x"a2",
         10348 => x"00",
         10349 => x"00",
         10350 => x"a2",
         10351 => x"00",
         10352 => x"00",
         10353 => x"a2",
         10354 => x"00",
         10355 => x"00",
         10356 => x"a2",
         10357 => x"00",
         10358 => x"00",
         10359 => x"a2",
         10360 => x"00",
         10361 => x"00",
         10362 => x"a2",
         10363 => x"00",
         10364 => x"00",
         10365 => x"a2",
         10366 => x"00",
         10367 => x"00",
         10368 => x"a2",
         10369 => x"00",
         10370 => x"00",
         10371 => x"a2",
         10372 => x"00",
         10373 => x"00",
         10374 => x"a2",
         10375 => x"00",
         10376 => x"00",
         10377 => x"a2",
         10378 => x"00",
         10379 => x"00",
         10380 => x"a2",
         10381 => x"00",
         10382 => x"00",
         10383 => x"a2",
         10384 => x"00",
         10385 => x"00",
         10386 => x"a2",
         10387 => x"00",
         10388 => x"00",
         10389 => x"a2",
         10390 => x"00",
         10391 => x"00",
         10392 => x"a2",
         10393 => x"00",
         10394 => x"00",
         10395 => x"a2",
         10396 => x"00",
         10397 => x"00",
         10398 => x"a2",
         10399 => x"00",
         10400 => x"00",
         10401 => x"a2",
         10402 => x"00",
         10403 => x"00",
         10404 => x"a2",
         10405 => x"00",
         10406 => x"00",
         10407 => x"44",
         10408 => x"43",
         10409 => x"42",
         10410 => x"41",
         10411 => x"36",
         10412 => x"35",
         10413 => x"34",
         10414 => x"46",
         10415 => x"33",
         10416 => x"32",
         10417 => x"31",
         10418 => x"00",
         10419 => x"00",
         10420 => x"00",
         10421 => x"00",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"73",
         10430 => x"79",
         10431 => x"73",
         10432 => x"00",
         10433 => x"00",
         10434 => x"34",
         10435 => x"20",
         10436 => x"00",
         10437 => x"69",
         10438 => x"20",
         10439 => x"72",
         10440 => x"74",
         10441 => x"65",
         10442 => x"73",
         10443 => x"79",
         10444 => x"6c",
         10445 => x"6f",
         10446 => x"46",
         10447 => x"00",
         10448 => x"6e",
         10449 => x"20",
         10450 => x"6e",
         10451 => x"65",
         10452 => x"20",
         10453 => x"74",
         10454 => x"20",
         10455 => x"65",
         10456 => x"69",
         10457 => x"6c",
         10458 => x"2e",
         10459 => x"00",
         10460 => x"3a",
         10461 => x"7c",
         10462 => x"00",
         10463 => x"3b",
         10464 => x"00",
         10465 => x"54",
         10466 => x"54",
         10467 => x"00",
         10468 => x"90",
         10469 => x"4f",
         10470 => x"30",
         10471 => x"20",
         10472 => x"45",
         10473 => x"20",
         10474 => x"33",
         10475 => x"20",
         10476 => x"20",
         10477 => x"45",
         10478 => x"20",
         10479 => x"20",
         10480 => x"20",
         10481 => x"a3",
         10482 => x"00",
         10483 => x"00",
         10484 => x"00",
         10485 => x"05",
         10486 => x"10",
         10487 => x"18",
         10488 => x"00",
         10489 => x"45",
         10490 => x"8f",
         10491 => x"45",
         10492 => x"8e",
         10493 => x"92",
         10494 => x"55",
         10495 => x"9a",
         10496 => x"9e",
         10497 => x"4f",
         10498 => x"a6",
         10499 => x"aa",
         10500 => x"ae",
         10501 => x"b2",
         10502 => x"b6",
         10503 => x"ba",
         10504 => x"be",
         10505 => x"c2",
         10506 => x"c6",
         10507 => x"ca",
         10508 => x"ce",
         10509 => x"d2",
         10510 => x"d6",
         10511 => x"da",
         10512 => x"de",
         10513 => x"e2",
         10514 => x"e6",
         10515 => x"ea",
         10516 => x"ee",
         10517 => x"f2",
         10518 => x"f6",
         10519 => x"fa",
         10520 => x"fe",
         10521 => x"2c",
         10522 => x"5d",
         10523 => x"2a",
         10524 => x"3f",
         10525 => x"00",
         10526 => x"00",
         10527 => x"00",
         10528 => x"02",
         10529 => x"00",
         10530 => x"00",
         10531 => x"00",
         10532 => x"00",
         10533 => x"00",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"00",
         10538 => x"00",
         10539 => x"00",
         10540 => x"00",
         10541 => x"00",
         10542 => x"00",
         10543 => x"00",
         10544 => x"00",
         10545 => x"00",
         10546 => x"00",
         10547 => x"00",
         10548 => x"00",
         10549 => x"01",
         10550 => x"00",
         10551 => x"00",
         10552 => x"00",
         10553 => x"00",
         10554 => x"23",
         10555 => x"00",
         10556 => x"00",
         10557 => x"00",
         10558 => x"25",
         10559 => x"25",
         10560 => x"25",
         10561 => x"25",
         10562 => x"25",
         10563 => x"25",
         10564 => x"25",
         10565 => x"25",
         10566 => x"25",
         10567 => x"25",
         10568 => x"25",
         10569 => x"25",
         10570 => x"25",
         10571 => x"25",
         10572 => x"25",
         10573 => x"25",
         10574 => x"25",
         10575 => x"25",
         10576 => x"25",
         10577 => x"25",
         10578 => x"25",
         10579 => x"25",
         10580 => x"25",
         10581 => x"25",
         10582 => x"00",
         10583 => x"03",
         10584 => x"03",
         10585 => x"03",
         10586 => x"03",
         10587 => x"03",
         10588 => x"03",
         10589 => x"22",
         10590 => x"00",
         10591 => x"22",
         10592 => x"23",
         10593 => x"22",
         10594 => x"22",
         10595 => x"22",
         10596 => x"00",
         10597 => x"00",
         10598 => x"03",
         10599 => x"03",
         10600 => x"03",
         10601 => x"00",
         10602 => x"01",
         10603 => x"01",
         10604 => x"01",
         10605 => x"01",
         10606 => x"01",
         10607 => x"01",
         10608 => x"02",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"01",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"02",
         10622 => x"01",
         10623 => x"02",
         10624 => x"01",
         10625 => x"01",
         10626 => x"01",
         10627 => x"01",
         10628 => x"01",
         10629 => x"01",
         10630 => x"01",
         10631 => x"01",
         10632 => x"01",
         10633 => x"01",
         10634 => x"01",
         10635 => x"01",
         10636 => x"01",
         10637 => x"01",
         10638 => x"01",
         10639 => x"01",
         10640 => x"01",
         10641 => x"01",
         10642 => x"01",
         10643 => x"01",
         10644 => x"01",
         10645 => x"01",
         10646 => x"01",
         10647 => x"01",
         10648 => x"00",
         10649 => x"01",
         10650 => x"01",
         10651 => x"01",
         10652 => x"01",
         10653 => x"01",
         10654 => x"01",
         10655 => x"00",
         10656 => x"02",
         10657 => x"02",
         10658 => x"02",
         10659 => x"02",
         10660 => x"02",
         10661 => x"02",
         10662 => x"01",
         10663 => x"02",
         10664 => x"01",
         10665 => x"01",
         10666 => x"01",
         10667 => x"02",
         10668 => x"02",
         10669 => x"02",
         10670 => x"01",
         10671 => x"02",
         10672 => x"02",
         10673 => x"01",
         10674 => x"2c",
         10675 => x"02",
         10676 => x"01",
         10677 => x"02",
         10678 => x"02",
         10679 => x"01",
         10680 => x"02",
         10681 => x"02",
         10682 => x"02",
         10683 => x"2c",
         10684 => x"02",
         10685 => x"02",
         10686 => x"01",
         10687 => x"02",
         10688 => x"02",
         10689 => x"02",
         10690 => x"01",
         10691 => x"02",
         10692 => x"02",
         10693 => x"02",
         10694 => x"03",
         10695 => x"03",
         10696 => x"03",
         10697 => x"00",
         10698 => x"03",
         10699 => x"03",
         10700 => x"03",
         10701 => x"00",
         10702 => x"03",
         10703 => x"03",
         10704 => x"00",
         10705 => x"03",
         10706 => x"03",
         10707 => x"03",
         10708 => x"03",
         10709 => x"03",
         10710 => x"03",
         10711 => x"03",
         10712 => x"03",
         10713 => x"04",
         10714 => x"04",
         10715 => x"04",
         10716 => x"04",
         10717 => x"04",
         10718 => x"04",
         10719 => x"04",
         10720 => x"01",
         10721 => x"04",
         10722 => x"00",
         10723 => x"00",
         10724 => x"1e",
         10725 => x"1e",
         10726 => x"1f",
         10727 => x"1f",
         10728 => x"1f",
         10729 => x"1f",
         10730 => x"1f",
         10731 => x"1f",
         10732 => x"1f",
         10733 => x"1f",
         10734 => x"1f",
         10735 => x"1f",
         10736 => x"06",
         10737 => x"00",
         10738 => x"1f",
         10739 => x"1f",
         10740 => x"1f",
         10741 => x"1f",
         10742 => x"1f",
         10743 => x"1f",
         10744 => x"1f",
         10745 => x"06",
         10746 => x"06",
         10747 => x"06",
         10748 => x"00",
         10749 => x"1f",
         10750 => x"1f",
         10751 => x"00",
         10752 => x"1f",
         10753 => x"1f",
         10754 => x"1f",
         10755 => x"1f",
         10756 => x"00",
         10757 => x"21",
         10758 => x"21",
         10759 => x"02",
         10760 => x"00",
         10761 => x"24",
         10762 => x"2c",
         10763 => x"2c",
         10764 => x"2c",
         10765 => x"2c",
         10766 => x"2c",
         10767 => x"2d",
         10768 => x"ff",
         10769 => x"00",
         10770 => x"00",
         10771 => x"98",
         10772 => x"01",
         10773 => x"00",
         10774 => x"00",
         10775 => x"98",
         10776 => x"01",
         10777 => x"00",
         10778 => x"00",
         10779 => x"98",
         10780 => x"03",
         10781 => x"00",
         10782 => x"00",
         10783 => x"98",
         10784 => x"03",
         10785 => x"00",
         10786 => x"00",
         10787 => x"98",
         10788 => x"03",
         10789 => x"00",
         10790 => x"00",
         10791 => x"98",
         10792 => x"04",
         10793 => x"00",
         10794 => x"00",
         10795 => x"98",
         10796 => x"04",
         10797 => x"00",
         10798 => x"00",
         10799 => x"98",
         10800 => x"04",
         10801 => x"00",
         10802 => x"00",
         10803 => x"98",
         10804 => x"04",
         10805 => x"00",
         10806 => x"00",
         10807 => x"98",
         10808 => x"04",
         10809 => x"00",
         10810 => x"00",
         10811 => x"98",
         10812 => x"04",
         10813 => x"00",
         10814 => x"00",
         10815 => x"98",
         10816 => x"04",
         10817 => x"00",
         10818 => x"00",
         10819 => x"98",
         10820 => x"05",
         10821 => x"00",
         10822 => x"00",
         10823 => x"98",
         10824 => x"05",
         10825 => x"00",
         10826 => x"00",
         10827 => x"98",
         10828 => x"05",
         10829 => x"00",
         10830 => x"00",
         10831 => x"99",
         10832 => x"05",
         10833 => x"00",
         10834 => x"00",
         10835 => x"99",
         10836 => x"07",
         10837 => x"00",
         10838 => x"00",
         10839 => x"99",
         10840 => x"07",
         10841 => x"00",
         10842 => x"00",
         10843 => x"99",
         10844 => x"08",
         10845 => x"00",
         10846 => x"00",
         10847 => x"99",
         10848 => x"08",
         10849 => x"00",
         10850 => x"00",
         10851 => x"99",
         10852 => x"08",
         10853 => x"00",
         10854 => x"00",
         10855 => x"99",
         10856 => x"08",
         10857 => x"00",
         10858 => x"00",
         10859 => x"99",
         10860 => x"09",
         10861 => x"00",
         10862 => x"00",
         10863 => x"99",
         10864 => x"09",
         10865 => x"00",
         10866 => x"00",
         10867 => x"99",
         10868 => x"09",
         10869 => x"00",
         10870 => x"00",
         10871 => x"99",
         10872 => x"09",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"7f",
         10878 => x"00",
         10879 => x"7f",
         10880 => x"00",
         10881 => x"7f",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"ff",
         10886 => x"00",
         10887 => x"00",
         10888 => x"78",
         10889 => x"00",
         10890 => x"e1",
         10891 => x"e1",
         10892 => x"e1",
         10893 => x"00",
         10894 => x"01",
         10895 => x"01",
         10896 => x"10",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"a2",
         10923 => x"00",
         10924 => x"a2",
         10925 => x"00",
         10926 => x"a3",
         10927 => x"00",
         10928 => x"f2",
         10929 => x"f6",
         10930 => x"fa",
         10931 => x"fe",
         10932 => x"c2",
         10933 => x"c6",
         10934 => x"e5",
         10935 => x"ef",
         10936 => x"62",
         10937 => x"66",
         10938 => x"6b",
         10939 => x"2e",
         10940 => x"22",
         10941 => x"26",
         10942 => x"4f",
         10943 => x"57",
         10944 => x"02",
         10945 => x"06",
         10946 => x"0a",
         10947 => x"0e",
         10948 => x"12",
         10949 => x"16",
         10950 => x"1a",
         10951 => x"be",
         10952 => x"82",
         10953 => x"86",
         10954 => x"8a",
         10955 => x"8e",
         10956 => x"92",
         10957 => x"96",
         10958 => x"9a",
         10959 => x"a5",
         10960 => x"00",
         10961 => x"00",
         10962 => x"00",
         10963 => x"00",
         10964 => x"00",
         10965 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"84",
           389 => x"82",
           390 => x"b3",
           391 => x"d6",
           392 => x"80",
           393 => x"d6",
           394 => x"e3",
           395 => x"e4",
           396 => x"90",
           397 => x"e4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"84",
           404 => x"82",
           405 => x"b1",
           406 => x"d6",
           407 => x"80",
           408 => x"d6",
           409 => x"d0",
           410 => x"d6",
           411 => x"80",
           412 => x"d6",
           413 => x"cb",
           414 => x"d6",
           415 => x"80",
           416 => x"d6",
           417 => x"d8",
           418 => x"e4",
           419 => x"90",
           420 => x"e4",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"84",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"84",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"84",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"84",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"84",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"84",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"84",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"84",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"84",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"84",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"84",
           467 => x"82",
           468 => x"82",
           469 => x"82",
           470 => x"84",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"84",
           475 => x"82",
           476 => x"82",
           477 => x"82",
           478 => x"84",
           479 => x"82",
           480 => x"82",
           481 => x"82",
           482 => x"84",
           483 => x"82",
           484 => x"82",
           485 => x"82",
           486 => x"84",
           487 => x"82",
           488 => x"82",
           489 => x"82",
           490 => x"84",
           491 => x"82",
           492 => x"82",
           493 => x"82",
           494 => x"84",
           495 => x"82",
           496 => x"82",
           497 => x"82",
           498 => x"84",
           499 => x"82",
           500 => x"82",
           501 => x"82",
           502 => x"84",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"84",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"84",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"84",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"84",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"84",
           523 => x"82",
           524 => x"82",
           525 => x"82",
           526 => x"84",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"84",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"84",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"84",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"84",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"84",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"84",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"84",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"84",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"84",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"84",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"84",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"84",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"84",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"84",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"84",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"84",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"84",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"84",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"ec",
           630 => x"d6",
           631 => x"82",
           632 => x"fb",
           633 => x"d6",
           634 => x"05",
           635 => x"e4",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"d8",
           644 => x"d6",
           645 => x"05",
           646 => x"e4",
           647 => x"08",
           648 => x"d8",
           649 => x"87",
           650 => x"d6",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"d6",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"e4",
           670 => x"0c",
           671 => x"d6",
           672 => x"05",
           673 => x"e4",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"e4",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"d6",
           696 => x"05",
           697 => x"e4",
           698 => x"08",
           699 => x"73",
           700 => x"e4",
           701 => x"08",
           702 => x"d6",
           703 => x"05",
           704 => x"e4",
           705 => x"08",
           706 => x"d6",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"d6",
           718 => x"3d",
           719 => x"e4",
           720 => x"d6",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"d6",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"d6",
           734 => x"05",
           735 => x"e4",
           736 => x"08",
           737 => x"e4",
           738 => x"08",
           739 => x"e4",
           740 => x"70",
           741 => x"81",
           742 => x"d6",
           743 => x"82",
           744 => x"dc",
           745 => x"d6",
           746 => x"05",
           747 => x"e4",
           748 => x"08",
           749 => x"80",
           750 => x"d6",
           751 => x"05",
           752 => x"d6",
           753 => x"8e",
           754 => x"d6",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"d6",
           761 => x"05",
           762 => x"e4",
           763 => x"08",
           764 => x"e4",
           765 => x"08",
           766 => x"e4",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"e4",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"e4",
           777 => x"d6",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"e4",
           797 => x"08",
           798 => x"53",
           799 => x"e4",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"e4",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"e4",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"d6",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"e4",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"d6",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"d6",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"d6",
           850 => x"05",
           851 => x"d6",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"e4",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"d6",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"e4",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"d6",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"d6",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"d6",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"d6",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"d6",
           943 => x"05",
           944 => x"51",
           945 => x"d6",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"d6",
           951 => x"05",
           952 => x"e4",
           953 => x"08",
           954 => x"d6",
           955 => x"05",
           956 => x"51",
           957 => x"d6",
           958 => x"05",
           959 => x"e4",
           960 => x"22",
           961 => x"53",
           962 => x"e4",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"d6",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"e4",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"d6",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"d6",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"d6",
          1003 => x"05",
          1004 => x"e4",
          1005 => x"08",
          1006 => x"d6",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"d6",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"e4",
          1025 => x"23",
          1026 => x"d6",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"d8",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"d6",
          1033 => x"05",
          1034 => x"d6",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"e4",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"d6",
          1046 => x"05",
          1047 => x"e4",
          1048 => x"08",
          1049 => x"d6",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"e4",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"e4",
          1059 => x"0c",
          1060 => x"d6",
          1061 => x"05",
          1062 => x"d6",
          1063 => x"05",
          1064 => x"e4",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"d6",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"e4",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"e4",
          1093 => x"34",
          1094 => x"d6",
          1095 => x"05",
          1096 => x"e4",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"d6",
          1102 => x"05",
          1103 => x"e4",
          1104 => x"08",
          1105 => x"d6",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"e4",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"e4",
          1115 => x"0c",
          1116 => x"d6",
          1117 => x"05",
          1118 => x"d6",
          1119 => x"05",
          1120 => x"e4",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"e4",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"d6",
          1132 => x"05",
          1133 => x"e4",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a5",
          1137 => x"d6",
          1138 => x"72",
          1139 => x"d6",
          1140 => x"05",
          1141 => x"e4",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"d6",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"d6",
          1160 => x"05",
          1161 => x"e4",
          1162 => x"08",
          1163 => x"e4",
          1164 => x"33",
          1165 => x"d6",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"d6",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"d6",
          1182 => x"05",
          1183 => x"e8",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"d6",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"d6",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"d6",
          1206 => x"05",
          1207 => x"e4",
          1208 => x"08",
          1209 => x"d6",
          1210 => x"05",
          1211 => x"e4",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"d6",
          1216 => x"05",
          1217 => x"53",
          1218 => x"e4",
          1219 => x"23",
          1220 => x"d6",
          1221 => x"05",
          1222 => x"53",
          1223 => x"e4",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"d6",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"e4",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"e4",
          1242 => x"22",
          1243 => x"51",
          1244 => x"d6",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"d6",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"d6",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"d6",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"d6",
          1287 => x"05",
          1288 => x"54",
          1289 => x"d6",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"d6",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"e4",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"d6",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"d6",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"d6",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"e4",
          1331 => x"08",
          1332 => x"89",
          1333 => x"d6",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"d6",
          1338 => x"05",
          1339 => x"d6",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"e4",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"d6",
          1348 => x"05",
          1349 => x"54",
          1350 => x"d6",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"d6",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"e4",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"d6",
          1365 => x"05",
          1366 => x"54",
          1367 => x"d6",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"d6",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"e4",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"d6",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"e4",
          1416 => x"08",
          1417 => x"e4",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"d6",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"e4",
          1439 => x"08",
          1440 => x"e4",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"d6",
          1449 => x"05",
          1450 => x"e8",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"e4",
          1468 => x"22",
          1469 => x"54",
          1470 => x"e4",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"e4",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"e4",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"e4",
          1492 => x"23",
          1493 => x"d6",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"d6",
          1501 => x"05",
          1502 => x"d6",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"d6",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"e4",
          1530 => x"d6",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"f2",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"d6",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"d6",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"bc",
          1556 => x"bc",
          1557 => x"d6",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"d8",
          1562 => x"80",
          1563 => x"38",
          1564 => x"d6",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"d6",
          1572 => x"72",
          1573 => x"38",
          1574 => x"d6",
          1575 => x"05",
          1576 => x"e4",
          1577 => x"08",
          1578 => x"e4",
          1579 => x"0c",
          1580 => x"e4",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"e4",
          1587 => x"0d",
          1588 => x"d6",
          1589 => x"05",
          1590 => x"e4",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"d6",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"e4",
          1606 => x"0c",
          1607 => x"d6",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"d6",
          1614 => x"05",
          1615 => x"d6",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"d8",
          1620 => x"80",
          1621 => x"38",
          1622 => x"d6",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"d6",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"d6",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"e4",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"e4",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"d6",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"d6",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"d6",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"e4",
          1683 => x"08",
          1684 => x"e4",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"e4",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"d6",
          1711 => x"3d",
          1712 => x"e4",
          1713 => x"d6",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"d6",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"e4",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"e4",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"d6",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"e4",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"e4",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"d6",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"d6",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"e4",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"d6",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"d6",
          1801 => x"05",
          1802 => x"52",
          1803 => x"e4",
          1804 => x"34",
          1805 => x"d6",
          1806 => x"05",
          1807 => x"52",
          1808 => x"e4",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"e4",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"d6",
          1827 => x"05",
          1828 => x"d8",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"e4",
          1832 => x"d6",
          1833 => x"3d",
          1834 => x"e4",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"d6",
          1840 => x"05",
          1841 => x"e4",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"e4",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"d6",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"d6",
          1858 => x"05",
          1859 => x"d6",
          1860 => x"05",
          1861 => x"e4",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"d6",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"d6",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"d6",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"d6",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"e4",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"d6",
          1917 => x"05",
          1918 => x"d6",
          1919 => x"85",
          1920 => x"d6",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"d6",
          1927 => x"05",
          1928 => x"e4",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"e4",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"e4",
          1950 => x"d6",
          1951 => x"3d",
          1952 => x"e4",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"e4",
          1959 => x"08",
          1960 => x"d6",
          1961 => x"05",
          1962 => x"e4",
          1963 => x"08",
          1964 => x"72",
          1965 => x"e4",
          1966 => x"08",
          1967 => x"d6",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"d6",
          1973 => x"05",
          1974 => x"d6",
          1975 => x"84",
          1976 => x"d6",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"d6",
          1983 => x"05",
          1984 => x"e4",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"d6",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"e4",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"e4",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"e4",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"d6",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"d6",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"e4",
          2043 => x"08",
          2044 => x"d6",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"d6",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"d6",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"d6",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"d6",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"d6",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"e4",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"e4",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"d6",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"8c",
          2099 => x"82",
          2100 => x"88",
          2101 => x"81",
          2102 => x"d6",
          2103 => x"82",
          2104 => x"f8",
          2105 => x"d6",
          2106 => x"05",
          2107 => x"70",
          2108 => x"80",
          2109 => x"82",
          2110 => x"70",
          2111 => x"08",
          2112 => x"54",
          2113 => x"08",
          2114 => x"8c",
          2115 => x"82",
          2116 => x"f4",
          2117 => x"39",
          2118 => x"08",
          2119 => x"82",
          2120 => x"f8",
          2121 => x"54",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"82",
          2125 => x"88",
          2126 => x"82",
          2127 => x"fc",
          2128 => x"fb",
          2129 => x"d6",
          2130 => x"82",
          2131 => x"f4",
          2132 => x"82",
          2133 => x"f4",
          2134 => x"d6",
          2135 => x"3d",
          2136 => x"e4",
          2137 => x"d6",
          2138 => x"82",
          2139 => x"fd",
          2140 => x"d6",
          2141 => x"05",
          2142 => x"e4",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"8d",
          2146 => x"82",
          2147 => x"fc",
          2148 => x"ec",
          2149 => x"e4",
          2150 => x"08",
          2151 => x"82",
          2152 => x"f8",
          2153 => x"05",
          2154 => x"08",
          2155 => x"70",
          2156 => x"51",
          2157 => x"2e",
          2158 => x"d6",
          2159 => x"05",
          2160 => x"82",
          2161 => x"8c",
          2162 => x"d6",
          2163 => x"05",
          2164 => x"84",
          2165 => x"39",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"e4",
          2169 => x"0c",
          2170 => x"08",
          2171 => x"82",
          2172 => x"88",
          2173 => x"70",
          2174 => x"08",
          2175 => x"51",
          2176 => x"08",
          2177 => x"82",
          2178 => x"85",
          2179 => x"d6",
          2180 => x"82",
          2181 => x"02",
          2182 => x"0c",
          2183 => x"82",
          2184 => x"88",
          2185 => x"d6",
          2186 => x"05",
          2187 => x"e4",
          2188 => x"08",
          2189 => x"d4",
          2190 => x"e4",
          2191 => x"08",
          2192 => x"d6",
          2193 => x"05",
          2194 => x"e4",
          2195 => x"08",
          2196 => x"d6",
          2197 => x"05",
          2198 => x"e4",
          2199 => x"08",
          2200 => x"38",
          2201 => x"08",
          2202 => x"51",
          2203 => x"e4",
          2204 => x"08",
          2205 => x"71",
          2206 => x"e4",
          2207 => x"08",
          2208 => x"d6",
          2209 => x"05",
          2210 => x"39",
          2211 => x"08",
          2212 => x"70",
          2213 => x"0c",
          2214 => x"0d",
          2215 => x"0c",
          2216 => x"e4",
          2217 => x"d6",
          2218 => x"3d",
          2219 => x"82",
          2220 => x"fc",
          2221 => x"d6",
          2222 => x"05",
          2223 => x"b9",
          2224 => x"e4",
          2225 => x"08",
          2226 => x"e4",
          2227 => x"0c",
          2228 => x"d6",
          2229 => x"05",
          2230 => x"e4",
          2231 => x"08",
          2232 => x"0b",
          2233 => x"08",
          2234 => x"82",
          2235 => x"f4",
          2236 => x"d6",
          2237 => x"05",
          2238 => x"e4",
          2239 => x"08",
          2240 => x"38",
          2241 => x"08",
          2242 => x"30",
          2243 => x"08",
          2244 => x"80",
          2245 => x"e4",
          2246 => x"0c",
          2247 => x"08",
          2248 => x"8a",
          2249 => x"82",
          2250 => x"f0",
          2251 => x"d6",
          2252 => x"05",
          2253 => x"e4",
          2254 => x"0c",
          2255 => x"d6",
          2256 => x"05",
          2257 => x"d6",
          2258 => x"05",
          2259 => x"c5",
          2260 => x"d8",
          2261 => x"d6",
          2262 => x"05",
          2263 => x"d6",
          2264 => x"05",
          2265 => x"90",
          2266 => x"e4",
          2267 => x"08",
          2268 => x"e4",
          2269 => x"0c",
          2270 => x"08",
          2271 => x"70",
          2272 => x"0c",
          2273 => x"0d",
          2274 => x"0c",
          2275 => x"e4",
          2276 => x"d6",
          2277 => x"3d",
          2278 => x"82",
          2279 => x"fc",
          2280 => x"d6",
          2281 => x"05",
          2282 => x"99",
          2283 => x"e4",
          2284 => x"08",
          2285 => x"e4",
          2286 => x"0c",
          2287 => x"d6",
          2288 => x"05",
          2289 => x"e4",
          2290 => x"08",
          2291 => x"38",
          2292 => x"08",
          2293 => x"30",
          2294 => x"08",
          2295 => x"81",
          2296 => x"e4",
          2297 => x"08",
          2298 => x"e4",
          2299 => x"08",
          2300 => x"3f",
          2301 => x"08",
          2302 => x"e4",
          2303 => x"0c",
          2304 => x"e4",
          2305 => x"08",
          2306 => x"38",
          2307 => x"08",
          2308 => x"30",
          2309 => x"08",
          2310 => x"82",
          2311 => x"f8",
          2312 => x"82",
          2313 => x"54",
          2314 => x"82",
          2315 => x"04",
          2316 => x"08",
          2317 => x"e4",
          2318 => x"0d",
          2319 => x"d6",
          2320 => x"05",
          2321 => x"d6",
          2322 => x"05",
          2323 => x"c5",
          2324 => x"d8",
          2325 => x"d6",
          2326 => x"85",
          2327 => x"d6",
          2328 => x"82",
          2329 => x"02",
          2330 => x"0c",
          2331 => x"81",
          2332 => x"e4",
          2333 => x"08",
          2334 => x"e4",
          2335 => x"08",
          2336 => x"82",
          2337 => x"70",
          2338 => x"0c",
          2339 => x"0d",
          2340 => x"0c",
          2341 => x"e4",
          2342 => x"d6",
          2343 => x"3d",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"0b",
          2347 => x"08",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"d6",
          2351 => x"05",
          2352 => x"38",
          2353 => x"08",
          2354 => x"80",
          2355 => x"80",
          2356 => x"e4",
          2357 => x"08",
          2358 => x"82",
          2359 => x"8c",
          2360 => x"82",
          2361 => x"8c",
          2362 => x"d6",
          2363 => x"05",
          2364 => x"d6",
          2365 => x"05",
          2366 => x"39",
          2367 => x"08",
          2368 => x"80",
          2369 => x"38",
          2370 => x"08",
          2371 => x"82",
          2372 => x"88",
          2373 => x"ad",
          2374 => x"e4",
          2375 => x"08",
          2376 => x"08",
          2377 => x"31",
          2378 => x"08",
          2379 => x"82",
          2380 => x"f8",
          2381 => x"d6",
          2382 => x"05",
          2383 => x"d6",
          2384 => x"05",
          2385 => x"e4",
          2386 => x"08",
          2387 => x"d6",
          2388 => x"05",
          2389 => x"e4",
          2390 => x"08",
          2391 => x"d6",
          2392 => x"05",
          2393 => x"39",
          2394 => x"08",
          2395 => x"80",
          2396 => x"82",
          2397 => x"88",
          2398 => x"82",
          2399 => x"f4",
          2400 => x"91",
          2401 => x"e4",
          2402 => x"08",
          2403 => x"e4",
          2404 => x"0c",
          2405 => x"e4",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"82",
          2409 => x"04",
          2410 => x"08",
          2411 => x"e4",
          2412 => x"0d",
          2413 => x"d6",
          2414 => x"05",
          2415 => x"e4",
          2416 => x"08",
          2417 => x"0c",
          2418 => x"08",
          2419 => x"70",
          2420 => x"72",
          2421 => x"82",
          2422 => x"f8",
          2423 => x"81",
          2424 => x"72",
          2425 => x"81",
          2426 => x"82",
          2427 => x"88",
          2428 => x"08",
          2429 => x"0c",
          2430 => x"82",
          2431 => x"f8",
          2432 => x"72",
          2433 => x"81",
          2434 => x"81",
          2435 => x"e4",
          2436 => x"34",
          2437 => x"08",
          2438 => x"70",
          2439 => x"71",
          2440 => x"51",
          2441 => x"82",
          2442 => x"f8",
          2443 => x"d6",
          2444 => x"05",
          2445 => x"b0",
          2446 => x"06",
          2447 => x"82",
          2448 => x"88",
          2449 => x"08",
          2450 => x"0c",
          2451 => x"53",
          2452 => x"d6",
          2453 => x"05",
          2454 => x"e4",
          2455 => x"33",
          2456 => x"08",
          2457 => x"82",
          2458 => x"e8",
          2459 => x"e2",
          2460 => x"82",
          2461 => x"e8",
          2462 => x"f8",
          2463 => x"80",
          2464 => x"0b",
          2465 => x"08",
          2466 => x"82",
          2467 => x"88",
          2468 => x"08",
          2469 => x"0c",
          2470 => x"53",
          2471 => x"d6",
          2472 => x"05",
          2473 => x"39",
          2474 => x"d6",
          2475 => x"05",
          2476 => x"e4",
          2477 => x"08",
          2478 => x"05",
          2479 => x"08",
          2480 => x"33",
          2481 => x"08",
          2482 => x"80",
          2483 => x"d6",
          2484 => x"05",
          2485 => x"a0",
          2486 => x"81",
          2487 => x"e4",
          2488 => x"0c",
          2489 => x"82",
          2490 => x"f8",
          2491 => x"af",
          2492 => x"38",
          2493 => x"08",
          2494 => x"53",
          2495 => x"83",
          2496 => x"80",
          2497 => x"e4",
          2498 => x"0c",
          2499 => x"88",
          2500 => x"e4",
          2501 => x"34",
          2502 => x"d6",
          2503 => x"05",
          2504 => x"73",
          2505 => x"82",
          2506 => x"f8",
          2507 => x"72",
          2508 => x"38",
          2509 => x"0b",
          2510 => x"08",
          2511 => x"82",
          2512 => x"0b",
          2513 => x"08",
          2514 => x"80",
          2515 => x"e4",
          2516 => x"0c",
          2517 => x"08",
          2518 => x"53",
          2519 => x"81",
          2520 => x"d6",
          2521 => x"05",
          2522 => x"e0",
          2523 => x"38",
          2524 => x"08",
          2525 => x"e0",
          2526 => x"72",
          2527 => x"08",
          2528 => x"82",
          2529 => x"f8",
          2530 => x"11",
          2531 => x"82",
          2532 => x"f8",
          2533 => x"d6",
          2534 => x"05",
          2535 => x"73",
          2536 => x"82",
          2537 => x"f8",
          2538 => x"11",
          2539 => x"82",
          2540 => x"f8",
          2541 => x"d6",
          2542 => x"05",
          2543 => x"89",
          2544 => x"80",
          2545 => x"e4",
          2546 => x"0c",
          2547 => x"82",
          2548 => x"f8",
          2549 => x"d6",
          2550 => x"05",
          2551 => x"72",
          2552 => x"38",
          2553 => x"d6",
          2554 => x"05",
          2555 => x"39",
          2556 => x"08",
          2557 => x"70",
          2558 => x"08",
          2559 => x"29",
          2560 => x"08",
          2561 => x"70",
          2562 => x"e4",
          2563 => x"0c",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"51",
          2568 => x"53",
          2569 => x"d6",
          2570 => x"05",
          2571 => x"39",
          2572 => x"08",
          2573 => x"53",
          2574 => x"90",
          2575 => x"e4",
          2576 => x"08",
          2577 => x"e4",
          2578 => x"0c",
          2579 => x"08",
          2580 => x"82",
          2581 => x"fc",
          2582 => x"0c",
          2583 => x"82",
          2584 => x"ec",
          2585 => x"d6",
          2586 => x"05",
          2587 => x"d8",
          2588 => x"0d",
          2589 => x"0c",
          2590 => x"e4",
          2591 => x"d6",
          2592 => x"3d",
          2593 => x"82",
          2594 => x"f0",
          2595 => x"d6",
          2596 => x"05",
          2597 => x"73",
          2598 => x"e4",
          2599 => x"08",
          2600 => x"53",
          2601 => x"72",
          2602 => x"08",
          2603 => x"72",
          2604 => x"53",
          2605 => x"09",
          2606 => x"38",
          2607 => x"08",
          2608 => x"70",
          2609 => x"71",
          2610 => x"39",
          2611 => x"08",
          2612 => x"53",
          2613 => x"09",
          2614 => x"38",
          2615 => x"d6",
          2616 => x"05",
          2617 => x"e4",
          2618 => x"08",
          2619 => x"05",
          2620 => x"08",
          2621 => x"33",
          2622 => x"08",
          2623 => x"82",
          2624 => x"f8",
          2625 => x"72",
          2626 => x"81",
          2627 => x"38",
          2628 => x"08",
          2629 => x"70",
          2630 => x"71",
          2631 => x"51",
          2632 => x"82",
          2633 => x"f8",
          2634 => x"d6",
          2635 => x"05",
          2636 => x"e4",
          2637 => x"0c",
          2638 => x"08",
          2639 => x"80",
          2640 => x"38",
          2641 => x"08",
          2642 => x"80",
          2643 => x"38",
          2644 => x"90",
          2645 => x"e4",
          2646 => x"34",
          2647 => x"08",
          2648 => x"70",
          2649 => x"71",
          2650 => x"51",
          2651 => x"82",
          2652 => x"f8",
          2653 => x"a4",
          2654 => x"82",
          2655 => x"f4",
          2656 => x"d6",
          2657 => x"05",
          2658 => x"81",
          2659 => x"70",
          2660 => x"72",
          2661 => x"e4",
          2662 => x"34",
          2663 => x"82",
          2664 => x"f8",
          2665 => x"72",
          2666 => x"38",
          2667 => x"d6",
          2668 => x"05",
          2669 => x"39",
          2670 => x"08",
          2671 => x"53",
          2672 => x"90",
          2673 => x"e4",
          2674 => x"33",
          2675 => x"26",
          2676 => x"39",
          2677 => x"d6",
          2678 => x"05",
          2679 => x"39",
          2680 => x"d6",
          2681 => x"05",
          2682 => x"82",
          2683 => x"f8",
          2684 => x"af",
          2685 => x"38",
          2686 => x"08",
          2687 => x"53",
          2688 => x"83",
          2689 => x"80",
          2690 => x"e4",
          2691 => x"0c",
          2692 => x"8a",
          2693 => x"e4",
          2694 => x"34",
          2695 => x"d6",
          2696 => x"05",
          2697 => x"e4",
          2698 => x"33",
          2699 => x"27",
          2700 => x"82",
          2701 => x"f8",
          2702 => x"80",
          2703 => x"94",
          2704 => x"e4",
          2705 => x"33",
          2706 => x"53",
          2707 => x"e4",
          2708 => x"34",
          2709 => x"08",
          2710 => x"d0",
          2711 => x"72",
          2712 => x"08",
          2713 => x"82",
          2714 => x"f8",
          2715 => x"90",
          2716 => x"38",
          2717 => x"08",
          2718 => x"f9",
          2719 => x"72",
          2720 => x"08",
          2721 => x"82",
          2722 => x"f8",
          2723 => x"72",
          2724 => x"38",
          2725 => x"d6",
          2726 => x"05",
          2727 => x"39",
          2728 => x"08",
          2729 => x"82",
          2730 => x"f4",
          2731 => x"54",
          2732 => x"8d",
          2733 => x"82",
          2734 => x"ec",
          2735 => x"f7",
          2736 => x"e4",
          2737 => x"33",
          2738 => x"e4",
          2739 => x"08",
          2740 => x"e4",
          2741 => x"33",
          2742 => x"d6",
          2743 => x"05",
          2744 => x"e4",
          2745 => x"08",
          2746 => x"05",
          2747 => x"08",
          2748 => x"55",
          2749 => x"82",
          2750 => x"f8",
          2751 => x"a5",
          2752 => x"e4",
          2753 => x"33",
          2754 => x"2e",
          2755 => x"d6",
          2756 => x"05",
          2757 => x"d6",
          2758 => x"05",
          2759 => x"e4",
          2760 => x"08",
          2761 => x"08",
          2762 => x"71",
          2763 => x"0b",
          2764 => x"08",
          2765 => x"82",
          2766 => x"ec",
          2767 => x"d6",
          2768 => x"3d",
          2769 => x"e4",
          2770 => x"3d",
          2771 => x"08",
          2772 => x"59",
          2773 => x"80",
          2774 => x"39",
          2775 => x"0c",
          2776 => x"54",
          2777 => x"74",
          2778 => x"a0",
          2779 => x"06",
          2780 => x"15",
          2781 => x"80",
          2782 => x"29",
          2783 => x"05",
          2784 => x"56",
          2785 => x"82",
          2786 => x"82",
          2787 => x"54",
          2788 => x"08",
          2789 => x"fc",
          2790 => x"d8",
          2791 => x"84",
          2792 => x"73",
          2793 => x"b4",
          2794 => x"70",
          2795 => x"58",
          2796 => x"27",
          2797 => x"54",
          2798 => x"d8",
          2799 => x"0d",
          2800 => x"0d",
          2801 => x"93",
          2802 => x"38",
          2803 => x"82",
          2804 => x"52",
          2805 => x"82",
          2806 => x"81",
          2807 => x"b2",
          2808 => x"f9",
          2809 => x"e8",
          2810 => x"39",
          2811 => x"51",
          2812 => x"82",
          2813 => x"80",
          2814 => x"b3",
          2815 => x"dd",
          2816 => x"ac",
          2817 => x"39",
          2818 => x"51",
          2819 => x"82",
          2820 => x"80",
          2821 => x"b3",
          2822 => x"c1",
          2823 => x"84",
          2824 => x"82",
          2825 => x"b5",
          2826 => x"b4",
          2827 => x"82",
          2828 => x"a9",
          2829 => x"ec",
          2830 => x"82",
          2831 => x"9d",
          2832 => x"9c",
          2833 => x"82",
          2834 => x"91",
          2835 => x"cc",
          2836 => x"82",
          2837 => x"85",
          2838 => x"f0",
          2839 => x"3f",
          2840 => x"04",
          2841 => x"77",
          2842 => x"74",
          2843 => x"8a",
          2844 => x"75",
          2845 => x"51",
          2846 => x"e8",
          2847 => x"ef",
          2848 => x"d6",
          2849 => x"75",
          2850 => x"3f",
          2851 => x"08",
          2852 => x"75",
          2853 => x"80",
          2854 => x"be",
          2855 => x"0d",
          2856 => x"0d",
          2857 => x"05",
          2858 => x"33",
          2859 => x"68",
          2860 => x"7a",
          2861 => x"51",
          2862 => x"78",
          2863 => x"ff",
          2864 => x"81",
          2865 => x"07",
          2866 => x"06",
          2867 => x"56",
          2868 => x"38",
          2869 => x"52",
          2870 => x"52",
          2871 => x"cf",
          2872 => x"d8",
          2873 => x"d6",
          2874 => x"38",
          2875 => x"08",
          2876 => x"88",
          2877 => x"d8",
          2878 => x"3d",
          2879 => x"84",
          2880 => x"52",
          2881 => x"97",
          2882 => x"d6",
          2883 => x"82",
          2884 => x"90",
          2885 => x"74",
          2886 => x"38",
          2887 => x"19",
          2888 => x"39",
          2889 => x"05",
          2890 => x"82",
          2891 => x"70",
          2892 => x"25",
          2893 => x"9f",
          2894 => x"51",
          2895 => x"74",
          2896 => x"38",
          2897 => x"53",
          2898 => x"88",
          2899 => x"51",
          2900 => x"76",
          2901 => x"d6",
          2902 => x"3d",
          2903 => x"3d",
          2904 => x"84",
          2905 => x"33",
          2906 => x"59",
          2907 => x"52",
          2908 => x"ad",
          2909 => x"d8",
          2910 => x"38",
          2911 => x"88",
          2912 => x"2e",
          2913 => x"39",
          2914 => x"57",
          2915 => x"56",
          2916 => x"55",
          2917 => x"08",
          2918 => x"bc",
          2919 => x"f2",
          2920 => x"82",
          2921 => x"ff",
          2922 => x"82",
          2923 => x"62",
          2924 => x"82",
          2925 => x"60",
          2926 => x"79",
          2927 => x"d8",
          2928 => x"39",
          2929 => x"82",
          2930 => x"8b",
          2931 => x"f3",
          2932 => x"61",
          2933 => x"05",
          2934 => x"33",
          2935 => x"68",
          2936 => x"5c",
          2937 => x"7a",
          2938 => x"e0",
          2939 => x"ea",
          2940 => x"e8",
          2941 => x"e2",
          2942 => x"74",
          2943 => x"80",
          2944 => x"2e",
          2945 => x"a0",
          2946 => x"80",
          2947 => x"18",
          2948 => x"27",
          2949 => x"22",
          2950 => x"ec",
          2951 => x"ba",
          2952 => x"82",
          2953 => x"ff",
          2954 => x"82",
          2955 => x"c3",
          2956 => x"53",
          2957 => x"8e",
          2958 => x"52",
          2959 => x"51",
          2960 => x"3f",
          2961 => x"b6",
          2962 => x"b7",
          2963 => x"15",
          2964 => x"74",
          2965 => x"7a",
          2966 => x"72",
          2967 => x"b7",
          2968 => x"b6",
          2969 => x"39",
          2970 => x"51",
          2971 => x"3f",
          2972 => x"82",
          2973 => x"52",
          2974 => x"b8",
          2975 => x"39",
          2976 => x"51",
          2977 => x"3f",
          2978 => x"79",
          2979 => x"38",
          2980 => x"33",
          2981 => x"56",
          2982 => x"83",
          2983 => x"80",
          2984 => x"27",
          2985 => x"53",
          2986 => x"70",
          2987 => x"51",
          2988 => x"2e",
          2989 => x"80",
          2990 => x"38",
          2991 => x"08",
          2992 => x"88",
          2993 => x"bc",
          2994 => x"51",
          2995 => x"81",
          2996 => x"b6",
          2997 => x"90",
          2998 => x"3f",
          2999 => x"1c",
          3000 => x"e7",
          3001 => x"d8",
          3002 => x"70",
          3003 => x"57",
          3004 => x"09",
          3005 => x"38",
          3006 => x"82",
          3007 => x"98",
          3008 => x"2c",
          3009 => x"70",
          3010 => x"32",
          3011 => x"72",
          3012 => x"07",
          3013 => x"58",
          3014 => x"57",
          3015 => x"d8",
          3016 => x"2e",
          3017 => x"85",
          3018 => x"8c",
          3019 => x"53",
          3020 => x"fd",
          3021 => x"53",
          3022 => x"d8",
          3023 => x"0d",
          3024 => x"0d",
          3025 => x"33",
          3026 => x"53",
          3027 => x"52",
          3028 => x"86",
          3029 => x"a4",
          3030 => x"c0",
          3031 => x"a4",
          3032 => x"b0",
          3033 => x"a5",
          3034 => x"b7",
          3035 => x"b4",
          3036 => x"80",
          3037 => x"a0",
          3038 => x"3d",
          3039 => x"3d",
          3040 => x"96",
          3041 => x"a5",
          3042 => x"51",
          3043 => x"82",
          3044 => x"99",
          3045 => x"51",
          3046 => x"72",
          3047 => x"81",
          3048 => x"71",
          3049 => x"38",
          3050 => x"9f",
          3051 => x"ec",
          3052 => x"3f",
          3053 => x"93",
          3054 => x"2a",
          3055 => x"51",
          3056 => x"2e",
          3057 => x"51",
          3058 => x"82",
          3059 => x"99",
          3060 => x"51",
          3061 => x"72",
          3062 => x"81",
          3063 => x"71",
          3064 => x"38",
          3065 => x"e3",
          3066 => x"8c",
          3067 => x"3f",
          3068 => x"d7",
          3069 => x"2a",
          3070 => x"51",
          3071 => x"2e",
          3072 => x"51",
          3073 => x"82",
          3074 => x"98",
          3075 => x"51",
          3076 => x"72",
          3077 => x"81",
          3078 => x"71",
          3079 => x"38",
          3080 => x"a7",
          3081 => x"b4",
          3082 => x"3f",
          3083 => x"9b",
          3084 => x"2a",
          3085 => x"51",
          3086 => x"2e",
          3087 => x"51",
          3088 => x"82",
          3089 => x"98",
          3090 => x"51",
          3091 => x"72",
          3092 => x"81",
          3093 => x"71",
          3094 => x"38",
          3095 => x"eb",
          3096 => x"dc",
          3097 => x"3f",
          3098 => x"df",
          3099 => x"2a",
          3100 => x"51",
          3101 => x"2e",
          3102 => x"51",
          3103 => x"82",
          3104 => x"97",
          3105 => x"51",
          3106 => x"a3",
          3107 => x"3d",
          3108 => x"3d",
          3109 => x"84",
          3110 => x"33",
          3111 => x"56",
          3112 => x"51",
          3113 => x"0b",
          3114 => x"c8",
          3115 => x"a9",
          3116 => x"82",
          3117 => x"82",
          3118 => x"81",
          3119 => x"82",
          3120 => x"30",
          3121 => x"d8",
          3122 => x"25",
          3123 => x"51",
          3124 => x"0b",
          3125 => x"c8",
          3126 => x"82",
          3127 => x"54",
          3128 => x"09",
          3129 => x"38",
          3130 => x"53",
          3131 => x"51",
          3132 => x"3f",
          3133 => x"08",
          3134 => x"38",
          3135 => x"08",
          3136 => x"3f",
          3137 => x"ed",
          3138 => x"97",
          3139 => x"0b",
          3140 => x"d0",
          3141 => x"0b",
          3142 => x"33",
          3143 => x"2e",
          3144 => x"8c",
          3145 => x"bc",
          3146 => x"75",
          3147 => x"3f",
          3148 => x"d6",
          3149 => x"3d",
          3150 => x"3d",
          3151 => x"41",
          3152 => x"82",
          3153 => x"5f",
          3154 => x"51",
          3155 => x"3f",
          3156 => x"08",
          3157 => x"59",
          3158 => x"09",
          3159 => x"38",
          3160 => x"83",
          3161 => x"c4",
          3162 => x"da",
          3163 => x"53",
          3164 => x"d8",
          3165 => x"88",
          3166 => x"d6",
          3167 => x"2e",
          3168 => x"b9",
          3169 => x"df",
          3170 => x"41",
          3171 => x"80",
          3172 => x"c6",
          3173 => x"70",
          3174 => x"f8",
          3175 => x"fd",
          3176 => x"3d",
          3177 => x"51",
          3178 => x"82",
          3179 => x"90",
          3180 => x"2c",
          3181 => x"80",
          3182 => x"a3",
          3183 => x"c2",
          3184 => x"78",
          3185 => x"d2",
          3186 => x"24",
          3187 => x"80",
          3188 => x"38",
          3189 => x"80",
          3190 => x"d6",
          3191 => x"c0",
          3192 => x"38",
          3193 => x"24",
          3194 => x"78",
          3195 => x"8c",
          3196 => x"39",
          3197 => x"2e",
          3198 => x"78",
          3199 => x"92",
          3200 => x"c3",
          3201 => x"38",
          3202 => x"2e",
          3203 => x"8a",
          3204 => x"81",
          3205 => x"88",
          3206 => x"83",
          3207 => x"78",
          3208 => x"89",
          3209 => x"8a",
          3210 => x"85",
          3211 => x"38",
          3212 => x"b5",
          3213 => x"11",
          3214 => x"05",
          3215 => x"3f",
          3216 => x"08",
          3217 => x"c5",
          3218 => x"fe",
          3219 => x"ff",
          3220 => x"ec",
          3221 => x"d6",
          3222 => x"2e",
          3223 => x"b5",
          3224 => x"11",
          3225 => x"05",
          3226 => x"3f",
          3227 => x"08",
          3228 => x"d6",
          3229 => x"82",
          3230 => x"ff",
          3231 => x"64",
          3232 => x"79",
          3233 => x"ec",
          3234 => x"78",
          3235 => x"05",
          3236 => x"7a",
          3237 => x"81",
          3238 => x"3d",
          3239 => x"53",
          3240 => x"51",
          3241 => x"82",
          3242 => x"80",
          3243 => x"38",
          3244 => x"fc",
          3245 => x"84",
          3246 => x"bd",
          3247 => x"d8",
          3248 => x"fd",
          3249 => x"3d",
          3250 => x"53",
          3251 => x"51",
          3252 => x"82",
          3253 => x"80",
          3254 => x"38",
          3255 => x"51",
          3256 => x"3f",
          3257 => x"64",
          3258 => x"38",
          3259 => x"70",
          3260 => x"33",
          3261 => x"81",
          3262 => x"39",
          3263 => x"80",
          3264 => x"84",
          3265 => x"f1",
          3266 => x"d8",
          3267 => x"fc",
          3268 => x"3d",
          3269 => x"53",
          3270 => x"51",
          3271 => x"82",
          3272 => x"80",
          3273 => x"38",
          3274 => x"f8",
          3275 => x"84",
          3276 => x"c5",
          3277 => x"d8",
          3278 => x"fc",
          3279 => x"ba",
          3280 => x"ad",
          3281 => x"5a",
          3282 => x"a8",
          3283 => x"33",
          3284 => x"5a",
          3285 => x"2e",
          3286 => x"55",
          3287 => x"33",
          3288 => x"82",
          3289 => x"ff",
          3290 => x"81",
          3291 => x"05",
          3292 => x"39",
          3293 => x"8f",
          3294 => x"39",
          3295 => x"80",
          3296 => x"84",
          3297 => x"f1",
          3298 => x"d8",
          3299 => x"38",
          3300 => x"33",
          3301 => x"2e",
          3302 => x"d3",
          3303 => x"80",
          3304 => x"d4",
          3305 => x"78",
          3306 => x"38",
          3307 => x"08",
          3308 => x"82",
          3309 => x"59",
          3310 => x"88",
          3311 => x"80",
          3312 => x"39",
          3313 => x"33",
          3314 => x"2e",
          3315 => x"d4",
          3316 => x"9a",
          3317 => x"b6",
          3318 => x"80",
          3319 => x"82",
          3320 => x"45",
          3321 => x"d4",
          3322 => x"80",
          3323 => x"3d",
          3324 => x"53",
          3325 => x"51",
          3326 => x"82",
          3327 => x"80",
          3328 => x"d4",
          3329 => x"78",
          3330 => x"38",
          3331 => x"08",
          3332 => x"39",
          3333 => x"33",
          3334 => x"2e",
          3335 => x"d3",
          3336 => x"bb",
          3337 => x"ba",
          3338 => x"80",
          3339 => x"82",
          3340 => x"44",
          3341 => x"d4",
          3342 => x"78",
          3343 => x"38",
          3344 => x"08",
          3345 => x"82",
          3346 => x"59",
          3347 => x"88",
          3348 => x"94",
          3349 => x"39",
          3350 => x"08",
          3351 => x"b5",
          3352 => x"11",
          3353 => x"05",
          3354 => x"3f",
          3355 => x"08",
          3356 => x"38",
          3357 => x"5c",
          3358 => x"83",
          3359 => x"7a",
          3360 => x"30",
          3361 => x"9f",
          3362 => x"06",
          3363 => x"5a",
          3364 => x"88",
          3365 => x"2e",
          3366 => x"43",
          3367 => x"51",
          3368 => x"a0",
          3369 => x"62",
          3370 => x"64",
          3371 => x"3f",
          3372 => x"51",
          3373 => x"b5",
          3374 => x"11",
          3375 => x"05",
          3376 => x"3f",
          3377 => x"08",
          3378 => x"c1",
          3379 => x"fe",
          3380 => x"ff",
          3381 => x"e7",
          3382 => x"d6",
          3383 => x"2e",
          3384 => x"59",
          3385 => x"05",
          3386 => x"64",
          3387 => x"b5",
          3388 => x"11",
          3389 => x"05",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"89",
          3393 => x"33",
          3394 => x"ba",
          3395 => x"a9",
          3396 => x"f2",
          3397 => x"80",
          3398 => x"51",
          3399 => x"3f",
          3400 => x"33",
          3401 => x"2e",
          3402 => x"9f",
          3403 => x"38",
          3404 => x"fc",
          3405 => x"84",
          3406 => x"bd",
          3407 => x"d8",
          3408 => x"91",
          3409 => x"02",
          3410 => x"33",
          3411 => x"81",
          3412 => x"b1",
          3413 => x"f0",
          3414 => x"3f",
          3415 => x"b5",
          3416 => x"11",
          3417 => x"05",
          3418 => x"3f",
          3419 => x"08",
          3420 => x"99",
          3421 => x"fe",
          3422 => x"ff",
          3423 => x"e0",
          3424 => x"d6",
          3425 => x"2e",
          3426 => x"59",
          3427 => x"05",
          3428 => x"82",
          3429 => x"78",
          3430 => x"fe",
          3431 => x"ff",
          3432 => x"e0",
          3433 => x"d6",
          3434 => x"38",
          3435 => x"61",
          3436 => x"52",
          3437 => x"51",
          3438 => x"3f",
          3439 => x"08",
          3440 => x"52",
          3441 => x"a8",
          3442 => x"46",
          3443 => x"78",
          3444 => x"b9",
          3445 => x"26",
          3446 => x"82",
          3447 => x"39",
          3448 => x"f0",
          3449 => x"84",
          3450 => x"bc",
          3451 => x"d8",
          3452 => x"93",
          3453 => x"02",
          3454 => x"22",
          3455 => x"05",
          3456 => x"42",
          3457 => x"82",
          3458 => x"c3",
          3459 => x"9f",
          3460 => x"fe",
          3461 => x"ff",
          3462 => x"df",
          3463 => x"d6",
          3464 => x"2e",
          3465 => x"b5",
          3466 => x"11",
          3467 => x"05",
          3468 => x"3f",
          3469 => x"08",
          3470 => x"38",
          3471 => x"0c",
          3472 => x"05",
          3473 => x"fe",
          3474 => x"ff",
          3475 => x"de",
          3476 => x"d6",
          3477 => x"38",
          3478 => x"61",
          3479 => x"52",
          3480 => x"51",
          3481 => x"3f",
          3482 => x"08",
          3483 => x"52",
          3484 => x"a7",
          3485 => x"46",
          3486 => x"78",
          3487 => x"8d",
          3488 => x"27",
          3489 => x"3d",
          3490 => x"53",
          3491 => x"51",
          3492 => x"82",
          3493 => x"80",
          3494 => x"61",
          3495 => x"59",
          3496 => x"42",
          3497 => x"82",
          3498 => x"c2",
          3499 => x"ab",
          3500 => x"ff",
          3501 => x"ff",
          3502 => x"e3",
          3503 => x"d6",
          3504 => x"2e",
          3505 => x"64",
          3506 => x"90",
          3507 => x"8a",
          3508 => x"78",
          3509 => x"ff",
          3510 => x"ff",
          3511 => x"e3",
          3512 => x"d6",
          3513 => x"2e",
          3514 => x"64",
          3515 => x"ac",
          3516 => x"e6",
          3517 => x"78",
          3518 => x"d8",
          3519 => x"f5",
          3520 => x"d6",
          3521 => x"82",
          3522 => x"ff",
          3523 => x"f4",
          3524 => x"bb",
          3525 => x"cd",
          3526 => x"9f",
          3527 => x"39",
          3528 => x"51",
          3529 => x"80",
          3530 => x"39",
          3531 => x"f4",
          3532 => x"3d",
          3533 => x"80",
          3534 => x"38",
          3535 => x"79",
          3536 => x"3f",
          3537 => x"08",
          3538 => x"d8",
          3539 => x"82",
          3540 => x"d6",
          3541 => x"b5",
          3542 => x"05",
          3543 => x"3f",
          3544 => x"08",
          3545 => x"5a",
          3546 => x"2e",
          3547 => x"82",
          3548 => x"51",
          3549 => x"82",
          3550 => x"8f",
          3551 => x"38",
          3552 => x"82",
          3553 => x"7a",
          3554 => x"38",
          3555 => x"8c",
          3556 => x"39",
          3557 => x"ad",
          3558 => x"39",
          3559 => x"56",
          3560 => x"bc",
          3561 => x"53",
          3562 => x"52",
          3563 => x"b0",
          3564 => x"a7",
          3565 => x"39",
          3566 => x"3d",
          3567 => x"51",
          3568 => x"ab",
          3569 => x"82",
          3570 => x"80",
          3571 => x"ac",
          3572 => x"ff",
          3573 => x"ff",
          3574 => x"93",
          3575 => x"80",
          3576 => x"b8",
          3577 => x"ff",
          3578 => x"ff",
          3579 => x"82",
          3580 => x"82",
          3581 => x"7c",
          3582 => x"80",
          3583 => x"80",
          3584 => x"80",
          3585 => x"ff",
          3586 => x"ea",
          3587 => x"d6",
          3588 => x"d6",
          3589 => x"70",
          3590 => x"07",
          3591 => x"5b",
          3592 => x"5a",
          3593 => x"83",
          3594 => x"78",
          3595 => x"78",
          3596 => x"38",
          3597 => x"81",
          3598 => x"59",
          3599 => x"38",
          3600 => x"7e",
          3601 => x"59",
          3602 => x"7e",
          3603 => x"81",
          3604 => x"82",
          3605 => x"ff",
          3606 => x"7c",
          3607 => x"3f",
          3608 => x"82",
          3609 => x"ff",
          3610 => x"f2",
          3611 => x"3d",
          3612 => x"82",
          3613 => x"87",
          3614 => x"08",
          3615 => x"80",
          3616 => x"d7",
          3617 => x"d6",
          3618 => x"2b",
          3619 => x"8c",
          3620 => x"87",
          3621 => x"73",
          3622 => x"3f",
          3623 => x"d8",
          3624 => x"c0",
          3625 => x"87",
          3626 => x"08",
          3627 => x"80",
          3628 => x"d6",
          3629 => x"d6",
          3630 => x"2b",
          3631 => x"9c",
          3632 => x"87",
          3633 => x"73",
          3634 => x"3f",
          3635 => x"d8",
          3636 => x"c0",
          3637 => x"8c",
          3638 => x"87",
          3639 => x"0c",
          3640 => x"0b",
          3641 => x"94",
          3642 => x"a0",
          3643 => x"73",
          3644 => x"55",
          3645 => x"af",
          3646 => x"f2",
          3647 => x"b0",
          3648 => x"8b",
          3649 => x"73",
          3650 => x"55",
          3651 => x"bf",
          3652 => x"ee",
          3653 => x"80",
          3654 => x"9e",
          3655 => x"80",
          3656 => x"96",
          3657 => x"80",
          3658 => x"8e",
          3659 => x"80",
          3660 => x"86",
          3661 => x"80",
          3662 => x"fe",
          3663 => x"8a",
          3664 => x"3f",
          3665 => x"51",
          3666 => x"81",
          3667 => x"81",
          3668 => x"83",
          3669 => x"95",
          3670 => x"5b",
          3671 => x"82",
          3672 => x"70",
          3673 => x"0c",
          3674 => x"0c",
          3675 => x"51",
          3676 => x"3f",
          3677 => x"91",
          3678 => x"bd",
          3679 => x"bc",
          3680 => x"bd",
          3681 => x"bc",
          3682 => x"de",
          3683 => x"d0",
          3684 => x"eb",
          3685 => x"a2",
          3686 => x"fe",
          3687 => x"52",
          3688 => x"88",
          3689 => x"d4",
          3690 => x"d8",
          3691 => x"06",
          3692 => x"14",
          3693 => x"80",
          3694 => x"71",
          3695 => x"0c",
          3696 => x"04",
          3697 => x"76",
          3698 => x"55",
          3699 => x"54",
          3700 => x"81",
          3701 => x"33",
          3702 => x"2e",
          3703 => x"86",
          3704 => x"53",
          3705 => x"33",
          3706 => x"2e",
          3707 => x"86",
          3708 => x"53",
          3709 => x"52",
          3710 => x"09",
          3711 => x"38",
          3712 => x"12",
          3713 => x"33",
          3714 => x"a2",
          3715 => x"81",
          3716 => x"2e",
          3717 => x"ea",
          3718 => x"81",
          3719 => x"72",
          3720 => x"70",
          3721 => x"38",
          3722 => x"80",
          3723 => x"73",
          3724 => x"72",
          3725 => x"70",
          3726 => x"81",
          3727 => x"81",
          3728 => x"32",
          3729 => x"80",
          3730 => x"51",
          3731 => x"80",
          3732 => x"80",
          3733 => x"05",
          3734 => x"75",
          3735 => x"70",
          3736 => x"0c",
          3737 => x"04",
          3738 => x"76",
          3739 => x"80",
          3740 => x"86",
          3741 => x"52",
          3742 => x"ac",
          3743 => x"d8",
          3744 => x"80",
          3745 => x"74",
          3746 => x"d6",
          3747 => x"3d",
          3748 => x"3d",
          3749 => x"11",
          3750 => x"52",
          3751 => x"70",
          3752 => x"98",
          3753 => x"33",
          3754 => x"82",
          3755 => x"26",
          3756 => x"84",
          3757 => x"83",
          3758 => x"26",
          3759 => x"85",
          3760 => x"84",
          3761 => x"26",
          3762 => x"86",
          3763 => x"85",
          3764 => x"26",
          3765 => x"88",
          3766 => x"86",
          3767 => x"e7",
          3768 => x"38",
          3769 => x"54",
          3770 => x"87",
          3771 => x"cc",
          3772 => x"87",
          3773 => x"0c",
          3774 => x"c0",
          3775 => x"82",
          3776 => x"c0",
          3777 => x"83",
          3778 => x"c0",
          3779 => x"84",
          3780 => x"c0",
          3781 => x"85",
          3782 => x"c0",
          3783 => x"86",
          3784 => x"c0",
          3785 => x"74",
          3786 => x"a4",
          3787 => x"c0",
          3788 => x"80",
          3789 => x"98",
          3790 => x"52",
          3791 => x"d8",
          3792 => x"0d",
          3793 => x"0d",
          3794 => x"c0",
          3795 => x"81",
          3796 => x"c0",
          3797 => x"5e",
          3798 => x"87",
          3799 => x"08",
          3800 => x"1c",
          3801 => x"98",
          3802 => x"79",
          3803 => x"87",
          3804 => x"08",
          3805 => x"1c",
          3806 => x"98",
          3807 => x"79",
          3808 => x"87",
          3809 => x"08",
          3810 => x"1c",
          3811 => x"98",
          3812 => x"7b",
          3813 => x"87",
          3814 => x"08",
          3815 => x"1c",
          3816 => x"0c",
          3817 => x"ff",
          3818 => x"83",
          3819 => x"58",
          3820 => x"57",
          3821 => x"56",
          3822 => x"55",
          3823 => x"54",
          3824 => x"53",
          3825 => x"ff",
          3826 => x"bd",
          3827 => x"9c",
          3828 => x"3d",
          3829 => x"3d",
          3830 => x"05",
          3831 => x"ec",
          3832 => x"ff",
          3833 => x"55",
          3834 => x"84",
          3835 => x"2e",
          3836 => x"c0",
          3837 => x"70",
          3838 => x"2a",
          3839 => x"53",
          3840 => x"80",
          3841 => x"71",
          3842 => x"81",
          3843 => x"70",
          3844 => x"81",
          3845 => x"06",
          3846 => x"80",
          3847 => x"71",
          3848 => x"81",
          3849 => x"70",
          3850 => x"73",
          3851 => x"51",
          3852 => x"80",
          3853 => x"2e",
          3854 => x"c0",
          3855 => x"74",
          3856 => x"82",
          3857 => x"87",
          3858 => x"ff",
          3859 => x"8f",
          3860 => x"30",
          3861 => x"51",
          3862 => x"82",
          3863 => x"83",
          3864 => x"f9",
          3865 => x"54",
          3866 => x"70",
          3867 => x"53",
          3868 => x"77",
          3869 => x"38",
          3870 => x"06",
          3871 => x"d3",
          3872 => x"81",
          3873 => x"57",
          3874 => x"c0",
          3875 => x"75",
          3876 => x"38",
          3877 => x"94",
          3878 => x"70",
          3879 => x"81",
          3880 => x"52",
          3881 => x"8c",
          3882 => x"2a",
          3883 => x"51",
          3884 => x"38",
          3885 => x"70",
          3886 => x"51",
          3887 => x"8d",
          3888 => x"2a",
          3889 => x"51",
          3890 => x"be",
          3891 => x"ff",
          3892 => x"c0",
          3893 => x"70",
          3894 => x"38",
          3895 => x"90",
          3896 => x"0c",
          3897 => x"33",
          3898 => x"06",
          3899 => x"70",
          3900 => x"76",
          3901 => x"0c",
          3902 => x"04",
          3903 => x"82",
          3904 => x"70",
          3905 => x"54",
          3906 => x"94",
          3907 => x"80",
          3908 => x"87",
          3909 => x"51",
          3910 => x"82",
          3911 => x"06",
          3912 => x"70",
          3913 => x"38",
          3914 => x"06",
          3915 => x"94",
          3916 => x"80",
          3917 => x"87",
          3918 => x"52",
          3919 => x"81",
          3920 => x"d6",
          3921 => x"84",
          3922 => x"fe",
          3923 => x"d3",
          3924 => x"81",
          3925 => x"53",
          3926 => x"84",
          3927 => x"2e",
          3928 => x"c0",
          3929 => x"71",
          3930 => x"2a",
          3931 => x"51",
          3932 => x"52",
          3933 => x"a0",
          3934 => x"ff",
          3935 => x"c0",
          3936 => x"70",
          3937 => x"38",
          3938 => x"90",
          3939 => x"70",
          3940 => x"98",
          3941 => x"51",
          3942 => x"d8",
          3943 => x"0d",
          3944 => x"0d",
          3945 => x"80",
          3946 => x"2a",
          3947 => x"51",
          3948 => x"84",
          3949 => x"c0",
          3950 => x"82",
          3951 => x"87",
          3952 => x"08",
          3953 => x"0c",
          3954 => x"94",
          3955 => x"f8",
          3956 => x"9e",
          3957 => x"d3",
          3958 => x"c0",
          3959 => x"82",
          3960 => x"87",
          3961 => x"08",
          3962 => x"0c",
          3963 => x"ac",
          3964 => x"88",
          3965 => x"9e",
          3966 => x"d4",
          3967 => x"c0",
          3968 => x"82",
          3969 => x"87",
          3970 => x"08",
          3971 => x"0c",
          3972 => x"bc",
          3973 => x"98",
          3974 => x"9e",
          3975 => x"d4",
          3976 => x"c0",
          3977 => x"82",
          3978 => x"87",
          3979 => x"08",
          3980 => x"d4",
          3981 => x"c0",
          3982 => x"82",
          3983 => x"87",
          3984 => x"08",
          3985 => x"0c",
          3986 => x"8c",
          3987 => x"b0",
          3988 => x"82",
          3989 => x"80",
          3990 => x"9e",
          3991 => x"84",
          3992 => x"51",
          3993 => x"80",
          3994 => x"81",
          3995 => x"d4",
          3996 => x"0b",
          3997 => x"90",
          3998 => x"80",
          3999 => x"52",
          4000 => x"2e",
          4001 => x"52",
          4002 => x"b6",
          4003 => x"87",
          4004 => x"08",
          4005 => x"0a",
          4006 => x"52",
          4007 => x"83",
          4008 => x"71",
          4009 => x"34",
          4010 => x"c0",
          4011 => x"70",
          4012 => x"06",
          4013 => x"70",
          4014 => x"38",
          4015 => x"82",
          4016 => x"80",
          4017 => x"9e",
          4018 => x"a0",
          4019 => x"51",
          4020 => x"80",
          4021 => x"81",
          4022 => x"d4",
          4023 => x"0b",
          4024 => x"90",
          4025 => x"80",
          4026 => x"52",
          4027 => x"2e",
          4028 => x"52",
          4029 => x"ba",
          4030 => x"87",
          4031 => x"08",
          4032 => x"80",
          4033 => x"52",
          4034 => x"83",
          4035 => x"71",
          4036 => x"34",
          4037 => x"c0",
          4038 => x"70",
          4039 => x"06",
          4040 => x"70",
          4041 => x"38",
          4042 => x"82",
          4043 => x"80",
          4044 => x"9e",
          4045 => x"81",
          4046 => x"51",
          4047 => x"80",
          4048 => x"81",
          4049 => x"d4",
          4050 => x"0b",
          4051 => x"90",
          4052 => x"c0",
          4053 => x"52",
          4054 => x"2e",
          4055 => x"52",
          4056 => x"be",
          4057 => x"87",
          4058 => x"08",
          4059 => x"06",
          4060 => x"70",
          4061 => x"38",
          4062 => x"82",
          4063 => x"87",
          4064 => x"08",
          4065 => x"06",
          4066 => x"51",
          4067 => x"82",
          4068 => x"80",
          4069 => x"9e",
          4070 => x"84",
          4071 => x"52",
          4072 => x"2e",
          4073 => x"52",
          4074 => x"c1",
          4075 => x"9e",
          4076 => x"83",
          4077 => x"84",
          4078 => x"51",
          4079 => x"c2",
          4080 => x"87",
          4081 => x"08",
          4082 => x"51",
          4083 => x"80",
          4084 => x"81",
          4085 => x"d4",
          4086 => x"c0",
          4087 => x"70",
          4088 => x"51",
          4089 => x"c4",
          4090 => x"0d",
          4091 => x"0d",
          4092 => x"51",
          4093 => x"3f",
          4094 => x"33",
          4095 => x"2e",
          4096 => x"bd",
          4097 => x"93",
          4098 => x"bd",
          4099 => x"af",
          4100 => x"d4",
          4101 => x"73",
          4102 => x"38",
          4103 => x"08",
          4104 => x"08",
          4105 => x"82",
          4106 => x"ff",
          4107 => x"82",
          4108 => x"54",
          4109 => x"94",
          4110 => x"88",
          4111 => x"8c",
          4112 => x"52",
          4113 => x"51",
          4114 => x"3f",
          4115 => x"33",
          4116 => x"2e",
          4117 => x"d3",
          4118 => x"d3",
          4119 => x"54",
          4120 => x"c0",
          4121 => x"f2",
          4122 => x"b9",
          4123 => x"80",
          4124 => x"82",
          4125 => x"82",
          4126 => x"11",
          4127 => x"be",
          4128 => x"92",
          4129 => x"d4",
          4130 => x"73",
          4131 => x"38",
          4132 => x"08",
          4133 => x"08",
          4134 => x"82",
          4135 => x"ff",
          4136 => x"82",
          4137 => x"54",
          4138 => x"8e",
          4139 => x"c0",
          4140 => x"bf",
          4141 => x"92",
          4142 => x"d4",
          4143 => x"73",
          4144 => x"38",
          4145 => x"33",
          4146 => x"b4",
          4147 => x"8a",
          4148 => x"c1",
          4149 => x"80",
          4150 => x"82",
          4151 => x"52",
          4152 => x"51",
          4153 => x"3f",
          4154 => x"33",
          4155 => x"2e",
          4156 => x"bf",
          4157 => x"ad",
          4158 => x"d4",
          4159 => x"73",
          4160 => x"38",
          4161 => x"51",
          4162 => x"3f",
          4163 => x"33",
          4164 => x"2e",
          4165 => x"c0",
          4166 => x"ad",
          4167 => x"d4",
          4168 => x"73",
          4169 => x"38",
          4170 => x"51",
          4171 => x"3f",
          4172 => x"33",
          4173 => x"2e",
          4174 => x"c0",
          4175 => x"ad",
          4176 => x"c0",
          4177 => x"ad",
          4178 => x"d4",
          4179 => x"82",
          4180 => x"ff",
          4181 => x"82",
          4182 => x"52",
          4183 => x"51",
          4184 => x"3f",
          4185 => x"08",
          4186 => x"8c",
          4187 => x"ea",
          4188 => x"b4",
          4189 => x"ed",
          4190 => x"a4",
          4191 => x"c1",
          4192 => x"90",
          4193 => x"d4",
          4194 => x"bd",
          4195 => x"75",
          4196 => x"3f",
          4197 => x"08",
          4198 => x"29",
          4199 => x"54",
          4200 => x"d8",
          4201 => x"c1",
          4202 => x"90",
          4203 => x"d4",
          4204 => x"73",
          4205 => x"38",
          4206 => x"08",
          4207 => x"c0",
          4208 => x"c4",
          4209 => x"d6",
          4210 => x"84",
          4211 => x"71",
          4212 => x"82",
          4213 => x"52",
          4214 => x"51",
          4215 => x"3f",
          4216 => x"33",
          4217 => x"2e",
          4218 => x"d4",
          4219 => x"bd",
          4220 => x"75",
          4221 => x"3f",
          4222 => x"08",
          4223 => x"29",
          4224 => x"54",
          4225 => x"d8",
          4226 => x"c2",
          4227 => x"8f",
          4228 => x"51",
          4229 => x"3f",
          4230 => x"04",
          4231 => x"02",
          4232 => x"ff",
          4233 => x"84",
          4234 => x"71",
          4235 => x"ad",
          4236 => x"71",
          4237 => x"c2",
          4238 => x"39",
          4239 => x"51",
          4240 => x"c2",
          4241 => x"39",
          4242 => x"51",
          4243 => x"c3",
          4244 => x"39",
          4245 => x"51",
          4246 => x"3f",
          4247 => x"04",
          4248 => x"0c",
          4249 => x"87",
          4250 => x"0c",
          4251 => x"c8",
          4252 => x"96",
          4253 => x"fd",
          4254 => x"98",
          4255 => x"2c",
          4256 => x"70",
          4257 => x"10",
          4258 => x"2b",
          4259 => x"54",
          4260 => x"0b",
          4261 => x"12",
          4262 => x"71",
          4263 => x"38",
          4264 => x"11",
          4265 => x"84",
          4266 => x"33",
          4267 => x"52",
          4268 => x"2e",
          4269 => x"83",
          4270 => x"72",
          4271 => x"0c",
          4272 => x"04",
          4273 => x"79",
          4274 => x"a3",
          4275 => x"33",
          4276 => x"72",
          4277 => x"38",
          4278 => x"08",
          4279 => x"ff",
          4280 => x"82",
          4281 => x"52",
          4282 => x"ad",
          4283 => x"f2",
          4284 => x"88",
          4285 => x"bc",
          4286 => x"ff",
          4287 => x"74",
          4288 => x"ff",
          4289 => x"39",
          4290 => x"8d",
          4291 => x"74",
          4292 => x"0d",
          4293 => x"0d",
          4294 => x"05",
          4295 => x"02",
          4296 => x"05",
          4297 => x"a4",
          4298 => x"29",
          4299 => x"05",
          4300 => x"59",
          4301 => x"59",
          4302 => x"86",
          4303 => x"9c",
          4304 => x"d5",
          4305 => x"84",
          4306 => x"cc",
          4307 => x"70",
          4308 => x"5a",
          4309 => x"82",
          4310 => x"75",
          4311 => x"a4",
          4312 => x"29",
          4313 => x"05",
          4314 => x"56",
          4315 => x"2e",
          4316 => x"53",
          4317 => x"51",
          4318 => x"3f",
          4319 => x"33",
          4320 => x"74",
          4321 => x"34",
          4322 => x"06",
          4323 => x"27",
          4324 => x"0b",
          4325 => x"34",
          4326 => x"b6",
          4327 => x"a0",
          4328 => x"80",
          4329 => x"82",
          4330 => x"55",
          4331 => x"8c",
          4332 => x"54",
          4333 => x"52",
          4334 => x"ec",
          4335 => x"d5",
          4336 => x"8a",
          4337 => x"80",
          4338 => x"a0",
          4339 => x"f0",
          4340 => x"3d",
          4341 => x"3d",
          4342 => x"cc",
          4343 => x"72",
          4344 => x"80",
          4345 => x"71",
          4346 => x"3f",
          4347 => x"ff",
          4348 => x"54",
          4349 => x"25",
          4350 => x"0b",
          4351 => x"34",
          4352 => x"08",
          4353 => x"2e",
          4354 => x"51",
          4355 => x"3f",
          4356 => x"08",
          4357 => x"3f",
          4358 => x"d5",
          4359 => x"3d",
          4360 => x"3d",
          4361 => x"80",
          4362 => x"a0",
          4363 => x"f6",
          4364 => x"d6",
          4365 => x"d3",
          4366 => x"a0",
          4367 => x"f8",
          4368 => x"70",
          4369 => x"9e",
          4370 => x"d6",
          4371 => x"2e",
          4372 => x"51",
          4373 => x"3f",
          4374 => x"08",
          4375 => x"82",
          4376 => x"25",
          4377 => x"d6",
          4378 => x"05",
          4379 => x"55",
          4380 => x"75",
          4381 => x"81",
          4382 => x"88",
          4383 => x"8a",
          4384 => x"ff",
          4385 => x"06",
          4386 => x"a6",
          4387 => x"d9",
          4388 => x"3d",
          4389 => x"08",
          4390 => x"70",
          4391 => x"52",
          4392 => x"08",
          4393 => x"c4",
          4394 => x"d8",
          4395 => x"38",
          4396 => x"d5",
          4397 => x"55",
          4398 => x"8b",
          4399 => x"56",
          4400 => x"3f",
          4401 => x"08",
          4402 => x"38",
          4403 => x"b2",
          4404 => x"d6",
          4405 => x"18",
          4406 => x"0b",
          4407 => x"08",
          4408 => x"82",
          4409 => x"ff",
          4410 => x"55",
          4411 => x"34",
          4412 => x"30",
          4413 => x"9f",
          4414 => x"55",
          4415 => x"85",
          4416 => x"ac",
          4417 => x"a0",
          4418 => x"08",
          4419 => x"f4",
          4420 => x"d6",
          4421 => x"2e",
          4422 => x"c6",
          4423 => x"89",
          4424 => x"77",
          4425 => x"06",
          4426 => x"52",
          4427 => x"b2",
          4428 => x"51",
          4429 => x"3f",
          4430 => x"54",
          4431 => x"08",
          4432 => x"58",
          4433 => x"d8",
          4434 => x"0d",
          4435 => x"0d",
          4436 => x"5c",
          4437 => x"57",
          4438 => x"73",
          4439 => x"81",
          4440 => x"78",
          4441 => x"56",
          4442 => x"98",
          4443 => x"70",
          4444 => x"33",
          4445 => x"73",
          4446 => x"81",
          4447 => x"75",
          4448 => x"38",
          4449 => x"88",
          4450 => x"a8",
          4451 => x"52",
          4452 => x"f3",
          4453 => x"d8",
          4454 => x"52",
          4455 => x"ff",
          4456 => x"82",
          4457 => x"80",
          4458 => x"15",
          4459 => x"81",
          4460 => x"74",
          4461 => x"38",
          4462 => x"e6",
          4463 => x"81",
          4464 => x"3d",
          4465 => x"f8",
          4466 => x"ad",
          4467 => x"d8",
          4468 => x"9a",
          4469 => x"53",
          4470 => x"51",
          4471 => x"82",
          4472 => x"81",
          4473 => x"74",
          4474 => x"54",
          4475 => x"14",
          4476 => x"06",
          4477 => x"74",
          4478 => x"38",
          4479 => x"82",
          4480 => x"8c",
          4481 => x"d3",
          4482 => x"3d",
          4483 => x"08",
          4484 => x"59",
          4485 => x"0b",
          4486 => x"82",
          4487 => x"82",
          4488 => x"55",
          4489 => x"cb",
          4490 => x"d5",
          4491 => x"55",
          4492 => x"81",
          4493 => x"2e",
          4494 => x"81",
          4495 => x"55",
          4496 => x"2e",
          4497 => x"a8",
          4498 => x"3f",
          4499 => x"08",
          4500 => x"0c",
          4501 => x"08",
          4502 => x"92",
          4503 => x"76",
          4504 => x"d8",
          4505 => x"df",
          4506 => x"d6",
          4507 => x"2e",
          4508 => x"c6",
          4509 => x"a2",
          4510 => x"f7",
          4511 => x"d8",
          4512 => x"d5",
          4513 => x"80",
          4514 => x"3d",
          4515 => x"81",
          4516 => x"82",
          4517 => x"56",
          4518 => x"08",
          4519 => x"81",
          4520 => x"38",
          4521 => x"08",
          4522 => x"db",
          4523 => x"d8",
          4524 => x"0b",
          4525 => x"08",
          4526 => x"82",
          4527 => x"ff",
          4528 => x"55",
          4529 => x"34",
          4530 => x"81",
          4531 => x"75",
          4532 => x"3f",
          4533 => x"81",
          4534 => x"54",
          4535 => x"83",
          4536 => x"74",
          4537 => x"81",
          4538 => x"38",
          4539 => x"82",
          4540 => x"76",
          4541 => x"d5",
          4542 => x"2e",
          4543 => x"d6",
          4544 => x"5d",
          4545 => x"82",
          4546 => x"98",
          4547 => x"2c",
          4548 => x"ff",
          4549 => x"78",
          4550 => x"82",
          4551 => x"70",
          4552 => x"98",
          4553 => x"90",
          4554 => x"2b",
          4555 => x"71",
          4556 => x"70",
          4557 => x"c3",
          4558 => x"08",
          4559 => x"51",
          4560 => x"59",
          4561 => x"5d",
          4562 => x"73",
          4563 => x"e9",
          4564 => x"27",
          4565 => x"81",
          4566 => x"81",
          4567 => x"70",
          4568 => x"55",
          4569 => x"80",
          4570 => x"53",
          4571 => x"51",
          4572 => x"82",
          4573 => x"81",
          4574 => x"73",
          4575 => x"38",
          4576 => x"90",
          4577 => x"b1",
          4578 => x"80",
          4579 => x"80",
          4580 => x"98",
          4581 => x"ff",
          4582 => x"55",
          4583 => x"97",
          4584 => x"74",
          4585 => x"f5",
          4586 => x"d6",
          4587 => x"ff",
          4588 => x"cc",
          4589 => x"80",
          4590 => x"2e",
          4591 => x"81",
          4592 => x"82",
          4593 => x"74",
          4594 => x"98",
          4595 => x"90",
          4596 => x"2b",
          4597 => x"70",
          4598 => x"82",
          4599 => x"98",
          4600 => x"51",
          4601 => x"58",
          4602 => x"77",
          4603 => x"06",
          4604 => x"82",
          4605 => x"08",
          4606 => x"0b",
          4607 => x"34",
          4608 => x"ee",
          4609 => x"39",
          4610 => x"94",
          4611 => x"ee",
          4612 => x"af",
          4613 => x"7d",
          4614 => x"73",
          4615 => x"e1",
          4616 => x"29",
          4617 => x"05",
          4618 => x"04",
          4619 => x"33",
          4620 => x"2e",
          4621 => x"82",
          4622 => x"55",
          4623 => x"ab",
          4624 => x"2b",
          4625 => x"51",
          4626 => x"24",
          4627 => x"1a",
          4628 => x"81",
          4629 => x"81",
          4630 => x"81",
          4631 => x"70",
          4632 => x"ee",
          4633 => x"51",
          4634 => x"82",
          4635 => x"81",
          4636 => x"74",
          4637 => x"34",
          4638 => x"ae",
          4639 => x"34",
          4640 => x"33",
          4641 => x"25",
          4642 => x"14",
          4643 => x"ee",
          4644 => x"ee",
          4645 => x"81",
          4646 => x"81",
          4647 => x"70",
          4648 => x"ee",
          4649 => x"51",
          4650 => x"77",
          4651 => x"82",
          4652 => x"52",
          4653 => x"33",
          4654 => x"a1",
          4655 => x"81",
          4656 => x"81",
          4657 => x"70",
          4658 => x"ee",
          4659 => x"51",
          4660 => x"24",
          4661 => x"ee",
          4662 => x"98",
          4663 => x"2c",
          4664 => x"33",
          4665 => x"56",
          4666 => x"fc",
          4667 => x"f2",
          4668 => x"88",
          4669 => x"bc",
          4670 => x"80",
          4671 => x"80",
          4672 => x"98",
          4673 => x"98",
          4674 => x"55",
          4675 => x"de",
          4676 => x"39",
          4677 => x"80",
          4678 => x"34",
          4679 => x"53",
          4680 => x"b6",
          4681 => x"9c",
          4682 => x"39",
          4683 => x"33",
          4684 => x"06",
          4685 => x"80",
          4686 => x"38",
          4687 => x"33",
          4688 => x"73",
          4689 => x"34",
          4690 => x"73",
          4691 => x"34",
          4692 => x"08",
          4693 => x"ff",
          4694 => x"82",
          4695 => x"70",
          4696 => x"98",
          4697 => x"98",
          4698 => x"56",
          4699 => x"25",
          4700 => x"1a",
          4701 => x"33",
          4702 => x"f2",
          4703 => x"73",
          4704 => x"a0",
          4705 => x"81",
          4706 => x"81",
          4707 => x"70",
          4708 => x"ee",
          4709 => x"51",
          4710 => x"24",
          4711 => x"f2",
          4712 => x"a0",
          4713 => x"8c",
          4714 => x"9c",
          4715 => x"2b",
          4716 => x"82",
          4717 => x"57",
          4718 => x"74",
          4719 => x"c1",
          4720 => x"bc",
          4721 => x"51",
          4722 => x"3f",
          4723 => x"0a",
          4724 => x"0a",
          4725 => x"2c",
          4726 => x"33",
          4727 => x"75",
          4728 => x"38",
          4729 => x"82",
          4730 => x"7a",
          4731 => x"74",
          4732 => x"bc",
          4733 => x"51",
          4734 => x"3f",
          4735 => x"52",
          4736 => x"c9",
          4737 => x"d8",
          4738 => x"06",
          4739 => x"38",
          4740 => x"33",
          4741 => x"2e",
          4742 => x"53",
          4743 => x"51",
          4744 => x"84",
          4745 => x"34",
          4746 => x"ee",
          4747 => x"0b",
          4748 => x"34",
          4749 => x"d8",
          4750 => x"0d",
          4751 => x"9c",
          4752 => x"80",
          4753 => x"38",
          4754 => x"08",
          4755 => x"ff",
          4756 => x"82",
          4757 => x"ff",
          4758 => x"82",
          4759 => x"73",
          4760 => x"54",
          4761 => x"ee",
          4762 => x"ee",
          4763 => x"55",
          4764 => x"f9",
          4765 => x"14",
          4766 => x"ee",
          4767 => x"98",
          4768 => x"2c",
          4769 => x"06",
          4770 => x"74",
          4771 => x"38",
          4772 => x"81",
          4773 => x"34",
          4774 => x"08",
          4775 => x"51",
          4776 => x"3f",
          4777 => x"0a",
          4778 => x"0a",
          4779 => x"2c",
          4780 => x"33",
          4781 => x"75",
          4782 => x"38",
          4783 => x"08",
          4784 => x"ff",
          4785 => x"82",
          4786 => x"70",
          4787 => x"98",
          4788 => x"98",
          4789 => x"56",
          4790 => x"24",
          4791 => x"82",
          4792 => x"52",
          4793 => x"9d",
          4794 => x"81",
          4795 => x"81",
          4796 => x"70",
          4797 => x"ee",
          4798 => x"51",
          4799 => x"25",
          4800 => x"fd",
          4801 => x"9c",
          4802 => x"ff",
          4803 => x"98",
          4804 => x"54",
          4805 => x"f7",
          4806 => x"f2",
          4807 => x"81",
          4808 => x"82",
          4809 => x"74",
          4810 => x"52",
          4811 => x"84",
          4812 => x"9c",
          4813 => x"ff",
          4814 => x"98",
          4815 => x"54",
          4816 => x"d6",
          4817 => x"39",
          4818 => x"53",
          4819 => x"b6",
          4820 => x"f0",
          4821 => x"82",
          4822 => x"80",
          4823 => x"98",
          4824 => x"39",
          4825 => x"82",
          4826 => x"55",
          4827 => x"a6",
          4828 => x"ff",
          4829 => x"82",
          4830 => x"82",
          4831 => x"82",
          4832 => x"81",
          4833 => x"05",
          4834 => x"79",
          4835 => x"d7",
          4836 => x"81",
          4837 => x"84",
          4838 => x"cc",
          4839 => x"08",
          4840 => x"80",
          4841 => x"74",
          4842 => x"db",
          4843 => x"d8",
          4844 => x"98",
          4845 => x"d8",
          4846 => x"06",
          4847 => x"74",
          4848 => x"ff",
          4849 => x"ff",
          4850 => x"fa",
          4851 => x"55",
          4852 => x"f6",
          4853 => x"51",
          4854 => x"3f",
          4855 => x"93",
          4856 => x"06",
          4857 => x"d4",
          4858 => x"74",
          4859 => x"38",
          4860 => x"a4",
          4861 => x"d6",
          4862 => x"ee",
          4863 => x"d6",
          4864 => x"ff",
          4865 => x"53",
          4866 => x"51",
          4867 => x"3f",
          4868 => x"7a",
          4869 => x"d4",
          4870 => x"08",
          4871 => x"80",
          4872 => x"74",
          4873 => x"df",
          4874 => x"d8",
          4875 => x"98",
          4876 => x"d8",
          4877 => x"06",
          4878 => x"74",
          4879 => x"ff",
          4880 => x"81",
          4881 => x"81",
          4882 => x"89",
          4883 => x"ee",
          4884 => x"7a",
          4885 => x"9c",
          4886 => x"98",
          4887 => x"51",
          4888 => x"f5",
          4889 => x"ee",
          4890 => x"81",
          4891 => x"ee",
          4892 => x"56",
          4893 => x"27",
          4894 => x"82",
          4895 => x"52",
          4896 => x"73",
          4897 => x"34",
          4898 => x"33",
          4899 => x"9a",
          4900 => x"ed",
          4901 => x"9c",
          4902 => x"80",
          4903 => x"38",
          4904 => x"08",
          4905 => x"ff",
          4906 => x"82",
          4907 => x"ff",
          4908 => x"82",
          4909 => x"f4",
          4910 => x"3d",
          4911 => x"05",
          4912 => x"8a",
          4913 => x"06",
          4914 => x"d6",
          4915 => x"05",
          4916 => x"0c",
          4917 => x"d6",
          4918 => x"87",
          4919 => x"82",
          4920 => x"80",
          4921 => x"c8",
          4922 => x"c4",
          4923 => x"82",
          4924 => x"05",
          4925 => x"82",
          4926 => x"05",
          4927 => x"80",
          4928 => x"d6",
          4929 => x"51",
          4930 => x"c0",
          4931 => x"34",
          4932 => x"08",
          4933 => x"d6",
          4934 => x"0b",
          4935 => x"08",
          4936 => x"82",
          4937 => x"81",
          4938 => x"c4",
          4939 => x"82",
          4940 => x"25",
          4941 => x"0b",
          4942 => x"0c",
          4943 => x"d6",
          4944 => x"0b",
          4945 => x"0c",
          4946 => x"04",
          4947 => x"d6",
          4948 => x"f9",
          4949 => x"bf",
          4950 => x"d6",
          4951 => x"80",
          4952 => x"cc",
          4953 => x"53",
          4954 => x"bf",
          4955 => x"a9",
          4956 => x"d6",
          4957 => x"80",
          4958 => x"34",
          4959 => x"81",
          4960 => x"d6",
          4961 => x"77",
          4962 => x"76",
          4963 => x"82",
          4964 => x"54",
          4965 => x"34",
          4966 => x"34",
          4967 => x"08",
          4968 => x"22",
          4969 => x"80",
          4970 => x"83",
          4971 => x"70",
          4972 => x"51",
          4973 => x"88",
          4974 => x"89",
          4975 => x"d6",
          4976 => x"88",
          4977 => x"d0",
          4978 => x"11",
          4979 => x"77",
          4980 => x"76",
          4981 => x"89",
          4982 => x"ff",
          4983 => x"52",
          4984 => x"72",
          4985 => x"fb",
          4986 => x"82",
          4987 => x"ff",
          4988 => x"51",
          4989 => x"d6",
          4990 => x"3d",
          4991 => x"3d",
          4992 => x"05",
          4993 => x"05",
          4994 => x"71",
          4995 => x"d0",
          4996 => x"2b",
          4997 => x"83",
          4998 => x"70",
          4999 => x"33",
          5000 => x"07",
          5001 => x"ae",
          5002 => x"81",
          5003 => x"07",
          5004 => x"53",
          5005 => x"54",
          5006 => x"53",
          5007 => x"77",
          5008 => x"18",
          5009 => x"d0",
          5010 => x"88",
          5011 => x"70",
          5012 => x"74",
          5013 => x"82",
          5014 => x"70",
          5015 => x"81",
          5016 => x"88",
          5017 => x"83",
          5018 => x"f8",
          5019 => x"56",
          5020 => x"73",
          5021 => x"06",
          5022 => x"54",
          5023 => x"82",
          5024 => x"81",
          5025 => x"72",
          5026 => x"82",
          5027 => x"16",
          5028 => x"34",
          5029 => x"34",
          5030 => x"04",
          5031 => x"82",
          5032 => x"02",
          5033 => x"05",
          5034 => x"2b",
          5035 => x"11",
          5036 => x"33",
          5037 => x"71",
          5038 => x"58",
          5039 => x"55",
          5040 => x"84",
          5041 => x"13",
          5042 => x"2b",
          5043 => x"2a",
          5044 => x"52",
          5045 => x"34",
          5046 => x"34",
          5047 => x"08",
          5048 => x"11",
          5049 => x"33",
          5050 => x"71",
          5051 => x"56",
          5052 => x"72",
          5053 => x"33",
          5054 => x"71",
          5055 => x"70",
          5056 => x"56",
          5057 => x"86",
          5058 => x"87",
          5059 => x"d6",
          5060 => x"70",
          5061 => x"33",
          5062 => x"07",
          5063 => x"ff",
          5064 => x"2a",
          5065 => x"53",
          5066 => x"34",
          5067 => x"34",
          5068 => x"04",
          5069 => x"02",
          5070 => x"82",
          5071 => x"71",
          5072 => x"11",
          5073 => x"12",
          5074 => x"2b",
          5075 => x"29",
          5076 => x"81",
          5077 => x"98",
          5078 => x"2b",
          5079 => x"53",
          5080 => x"56",
          5081 => x"71",
          5082 => x"f6",
          5083 => x"fe",
          5084 => x"d6",
          5085 => x"16",
          5086 => x"12",
          5087 => x"2b",
          5088 => x"07",
          5089 => x"33",
          5090 => x"71",
          5091 => x"70",
          5092 => x"ff",
          5093 => x"52",
          5094 => x"5a",
          5095 => x"05",
          5096 => x"54",
          5097 => x"13",
          5098 => x"13",
          5099 => x"d0",
          5100 => x"70",
          5101 => x"33",
          5102 => x"71",
          5103 => x"56",
          5104 => x"72",
          5105 => x"81",
          5106 => x"88",
          5107 => x"81",
          5108 => x"70",
          5109 => x"51",
          5110 => x"72",
          5111 => x"81",
          5112 => x"3d",
          5113 => x"3d",
          5114 => x"d0",
          5115 => x"05",
          5116 => x"70",
          5117 => x"11",
          5118 => x"83",
          5119 => x"8b",
          5120 => x"2b",
          5121 => x"59",
          5122 => x"73",
          5123 => x"81",
          5124 => x"88",
          5125 => x"8c",
          5126 => x"22",
          5127 => x"88",
          5128 => x"53",
          5129 => x"73",
          5130 => x"14",
          5131 => x"d0",
          5132 => x"70",
          5133 => x"33",
          5134 => x"71",
          5135 => x"56",
          5136 => x"72",
          5137 => x"33",
          5138 => x"71",
          5139 => x"70",
          5140 => x"55",
          5141 => x"82",
          5142 => x"83",
          5143 => x"d6",
          5144 => x"82",
          5145 => x"12",
          5146 => x"2b",
          5147 => x"d8",
          5148 => x"87",
          5149 => x"f7",
          5150 => x"82",
          5151 => x"31",
          5152 => x"83",
          5153 => x"70",
          5154 => x"fd",
          5155 => x"d6",
          5156 => x"83",
          5157 => x"82",
          5158 => x"12",
          5159 => x"2b",
          5160 => x"07",
          5161 => x"33",
          5162 => x"71",
          5163 => x"90",
          5164 => x"42",
          5165 => x"5b",
          5166 => x"54",
          5167 => x"8d",
          5168 => x"80",
          5169 => x"fe",
          5170 => x"84",
          5171 => x"33",
          5172 => x"71",
          5173 => x"83",
          5174 => x"11",
          5175 => x"53",
          5176 => x"55",
          5177 => x"34",
          5178 => x"06",
          5179 => x"14",
          5180 => x"d0",
          5181 => x"84",
          5182 => x"13",
          5183 => x"2b",
          5184 => x"2a",
          5185 => x"56",
          5186 => x"16",
          5187 => x"16",
          5188 => x"d0",
          5189 => x"80",
          5190 => x"34",
          5191 => x"14",
          5192 => x"d0",
          5193 => x"84",
          5194 => x"85",
          5195 => x"d6",
          5196 => x"70",
          5197 => x"33",
          5198 => x"07",
          5199 => x"80",
          5200 => x"2a",
          5201 => x"56",
          5202 => x"34",
          5203 => x"34",
          5204 => x"04",
          5205 => x"73",
          5206 => x"d0",
          5207 => x"f7",
          5208 => x"80",
          5209 => x"71",
          5210 => x"3f",
          5211 => x"04",
          5212 => x"80",
          5213 => x"f8",
          5214 => x"d6",
          5215 => x"ff",
          5216 => x"d6",
          5217 => x"11",
          5218 => x"33",
          5219 => x"07",
          5220 => x"56",
          5221 => x"ff",
          5222 => x"78",
          5223 => x"38",
          5224 => x"17",
          5225 => x"12",
          5226 => x"2b",
          5227 => x"ff",
          5228 => x"31",
          5229 => x"ff",
          5230 => x"27",
          5231 => x"56",
          5232 => x"79",
          5233 => x"73",
          5234 => x"38",
          5235 => x"5b",
          5236 => x"85",
          5237 => x"88",
          5238 => x"54",
          5239 => x"78",
          5240 => x"2e",
          5241 => x"79",
          5242 => x"76",
          5243 => x"d6",
          5244 => x"70",
          5245 => x"33",
          5246 => x"07",
          5247 => x"ff",
          5248 => x"5a",
          5249 => x"73",
          5250 => x"38",
          5251 => x"54",
          5252 => x"81",
          5253 => x"54",
          5254 => x"81",
          5255 => x"7a",
          5256 => x"06",
          5257 => x"51",
          5258 => x"81",
          5259 => x"80",
          5260 => x"52",
          5261 => x"c6",
          5262 => x"d0",
          5263 => x"86",
          5264 => x"12",
          5265 => x"2b",
          5266 => x"07",
          5267 => x"55",
          5268 => x"17",
          5269 => x"ff",
          5270 => x"2a",
          5271 => x"54",
          5272 => x"34",
          5273 => x"06",
          5274 => x"15",
          5275 => x"d0",
          5276 => x"2b",
          5277 => x"1e",
          5278 => x"87",
          5279 => x"88",
          5280 => x"88",
          5281 => x"5e",
          5282 => x"54",
          5283 => x"34",
          5284 => x"34",
          5285 => x"08",
          5286 => x"11",
          5287 => x"33",
          5288 => x"71",
          5289 => x"53",
          5290 => x"74",
          5291 => x"86",
          5292 => x"87",
          5293 => x"d6",
          5294 => x"16",
          5295 => x"11",
          5296 => x"33",
          5297 => x"07",
          5298 => x"53",
          5299 => x"56",
          5300 => x"16",
          5301 => x"16",
          5302 => x"d0",
          5303 => x"05",
          5304 => x"d6",
          5305 => x"3d",
          5306 => x"3d",
          5307 => x"82",
          5308 => x"84",
          5309 => x"3f",
          5310 => x"80",
          5311 => x"71",
          5312 => x"3f",
          5313 => x"08",
          5314 => x"d6",
          5315 => x"3d",
          5316 => x"3d",
          5317 => x"40",
          5318 => x"42",
          5319 => x"d0",
          5320 => x"09",
          5321 => x"38",
          5322 => x"7b",
          5323 => x"51",
          5324 => x"82",
          5325 => x"54",
          5326 => x"7e",
          5327 => x"51",
          5328 => x"7e",
          5329 => x"39",
          5330 => x"8f",
          5331 => x"d8",
          5332 => x"ff",
          5333 => x"d0",
          5334 => x"31",
          5335 => x"83",
          5336 => x"70",
          5337 => x"11",
          5338 => x"12",
          5339 => x"2b",
          5340 => x"31",
          5341 => x"ff",
          5342 => x"29",
          5343 => x"88",
          5344 => x"33",
          5345 => x"71",
          5346 => x"70",
          5347 => x"44",
          5348 => x"41",
          5349 => x"5b",
          5350 => x"5b",
          5351 => x"25",
          5352 => x"81",
          5353 => x"75",
          5354 => x"ff",
          5355 => x"54",
          5356 => x"83",
          5357 => x"88",
          5358 => x"88",
          5359 => x"33",
          5360 => x"71",
          5361 => x"90",
          5362 => x"47",
          5363 => x"54",
          5364 => x"8b",
          5365 => x"31",
          5366 => x"ff",
          5367 => x"77",
          5368 => x"fe",
          5369 => x"54",
          5370 => x"09",
          5371 => x"38",
          5372 => x"c0",
          5373 => x"ff",
          5374 => x"81",
          5375 => x"8e",
          5376 => x"24",
          5377 => x"51",
          5378 => x"81",
          5379 => x"18",
          5380 => x"24",
          5381 => x"79",
          5382 => x"33",
          5383 => x"71",
          5384 => x"53",
          5385 => x"f4",
          5386 => x"78",
          5387 => x"3f",
          5388 => x"08",
          5389 => x"06",
          5390 => x"53",
          5391 => x"82",
          5392 => x"11",
          5393 => x"55",
          5394 => x"d1",
          5395 => x"d0",
          5396 => x"05",
          5397 => x"ff",
          5398 => x"81",
          5399 => x"15",
          5400 => x"24",
          5401 => x"78",
          5402 => x"3f",
          5403 => x"08",
          5404 => x"33",
          5405 => x"71",
          5406 => x"53",
          5407 => x"9c",
          5408 => x"78",
          5409 => x"3f",
          5410 => x"08",
          5411 => x"06",
          5412 => x"53",
          5413 => x"82",
          5414 => x"11",
          5415 => x"55",
          5416 => x"f9",
          5417 => x"d0",
          5418 => x"05",
          5419 => x"19",
          5420 => x"83",
          5421 => x"58",
          5422 => x"7f",
          5423 => x"b0",
          5424 => x"d8",
          5425 => x"d6",
          5426 => x"2e",
          5427 => x"53",
          5428 => x"d6",
          5429 => x"ff",
          5430 => x"73",
          5431 => x"3f",
          5432 => x"78",
          5433 => x"80",
          5434 => x"78",
          5435 => x"3f",
          5436 => x"2b",
          5437 => x"08",
          5438 => x"51",
          5439 => x"7b",
          5440 => x"d6",
          5441 => x"3d",
          5442 => x"3d",
          5443 => x"29",
          5444 => x"fb",
          5445 => x"d6",
          5446 => x"82",
          5447 => x"80",
          5448 => x"73",
          5449 => x"82",
          5450 => x"51",
          5451 => x"3f",
          5452 => x"d8",
          5453 => x"0d",
          5454 => x"0d",
          5455 => x"33",
          5456 => x"70",
          5457 => x"38",
          5458 => x"11",
          5459 => x"82",
          5460 => x"83",
          5461 => x"fc",
          5462 => x"9b",
          5463 => x"84",
          5464 => x"33",
          5465 => x"51",
          5466 => x"80",
          5467 => x"84",
          5468 => x"92",
          5469 => x"51",
          5470 => x"80",
          5471 => x"81",
          5472 => x"72",
          5473 => x"92",
          5474 => x"81",
          5475 => x"0b",
          5476 => x"8c",
          5477 => x"71",
          5478 => x"06",
          5479 => x"80",
          5480 => x"87",
          5481 => x"08",
          5482 => x"38",
          5483 => x"80",
          5484 => x"71",
          5485 => x"c0",
          5486 => x"51",
          5487 => x"87",
          5488 => x"d6",
          5489 => x"82",
          5490 => x"33",
          5491 => x"d6",
          5492 => x"3d",
          5493 => x"3d",
          5494 => x"64",
          5495 => x"bf",
          5496 => x"40",
          5497 => x"74",
          5498 => x"cd",
          5499 => x"d8",
          5500 => x"7a",
          5501 => x"81",
          5502 => x"72",
          5503 => x"87",
          5504 => x"11",
          5505 => x"8c",
          5506 => x"92",
          5507 => x"5a",
          5508 => x"58",
          5509 => x"c0",
          5510 => x"76",
          5511 => x"76",
          5512 => x"70",
          5513 => x"81",
          5514 => x"54",
          5515 => x"8e",
          5516 => x"52",
          5517 => x"81",
          5518 => x"81",
          5519 => x"74",
          5520 => x"53",
          5521 => x"83",
          5522 => x"78",
          5523 => x"8f",
          5524 => x"2e",
          5525 => x"c0",
          5526 => x"52",
          5527 => x"87",
          5528 => x"08",
          5529 => x"2e",
          5530 => x"84",
          5531 => x"38",
          5532 => x"87",
          5533 => x"15",
          5534 => x"70",
          5535 => x"52",
          5536 => x"ff",
          5537 => x"39",
          5538 => x"81",
          5539 => x"ff",
          5540 => x"57",
          5541 => x"90",
          5542 => x"80",
          5543 => x"71",
          5544 => x"78",
          5545 => x"38",
          5546 => x"80",
          5547 => x"80",
          5548 => x"81",
          5549 => x"72",
          5550 => x"0c",
          5551 => x"04",
          5552 => x"60",
          5553 => x"8c",
          5554 => x"33",
          5555 => x"5b",
          5556 => x"74",
          5557 => x"e1",
          5558 => x"d8",
          5559 => x"79",
          5560 => x"78",
          5561 => x"06",
          5562 => x"77",
          5563 => x"87",
          5564 => x"11",
          5565 => x"8c",
          5566 => x"92",
          5567 => x"59",
          5568 => x"85",
          5569 => x"98",
          5570 => x"7d",
          5571 => x"0c",
          5572 => x"08",
          5573 => x"70",
          5574 => x"53",
          5575 => x"2e",
          5576 => x"70",
          5577 => x"33",
          5578 => x"18",
          5579 => x"2a",
          5580 => x"51",
          5581 => x"2e",
          5582 => x"c0",
          5583 => x"52",
          5584 => x"87",
          5585 => x"08",
          5586 => x"2e",
          5587 => x"84",
          5588 => x"38",
          5589 => x"87",
          5590 => x"15",
          5591 => x"70",
          5592 => x"52",
          5593 => x"ff",
          5594 => x"39",
          5595 => x"81",
          5596 => x"80",
          5597 => x"52",
          5598 => x"90",
          5599 => x"80",
          5600 => x"71",
          5601 => x"7a",
          5602 => x"38",
          5603 => x"80",
          5604 => x"80",
          5605 => x"81",
          5606 => x"72",
          5607 => x"0c",
          5608 => x"04",
          5609 => x"7a",
          5610 => x"a3",
          5611 => x"88",
          5612 => x"33",
          5613 => x"56",
          5614 => x"3f",
          5615 => x"08",
          5616 => x"83",
          5617 => x"fe",
          5618 => x"87",
          5619 => x"0c",
          5620 => x"76",
          5621 => x"38",
          5622 => x"93",
          5623 => x"2b",
          5624 => x"8c",
          5625 => x"71",
          5626 => x"38",
          5627 => x"71",
          5628 => x"c6",
          5629 => x"39",
          5630 => x"81",
          5631 => x"06",
          5632 => x"71",
          5633 => x"38",
          5634 => x"8c",
          5635 => x"e8",
          5636 => x"98",
          5637 => x"71",
          5638 => x"73",
          5639 => x"92",
          5640 => x"72",
          5641 => x"06",
          5642 => x"f7",
          5643 => x"80",
          5644 => x"88",
          5645 => x"0c",
          5646 => x"80",
          5647 => x"56",
          5648 => x"56",
          5649 => x"82",
          5650 => x"88",
          5651 => x"fe",
          5652 => x"81",
          5653 => x"33",
          5654 => x"07",
          5655 => x"0c",
          5656 => x"3d",
          5657 => x"3d",
          5658 => x"11",
          5659 => x"33",
          5660 => x"71",
          5661 => x"81",
          5662 => x"72",
          5663 => x"75",
          5664 => x"82",
          5665 => x"52",
          5666 => x"54",
          5667 => x"0d",
          5668 => x"0d",
          5669 => x"05",
          5670 => x"52",
          5671 => x"70",
          5672 => x"34",
          5673 => x"51",
          5674 => x"83",
          5675 => x"ff",
          5676 => x"75",
          5677 => x"72",
          5678 => x"54",
          5679 => x"2a",
          5680 => x"70",
          5681 => x"34",
          5682 => x"51",
          5683 => x"81",
          5684 => x"70",
          5685 => x"70",
          5686 => x"3d",
          5687 => x"3d",
          5688 => x"77",
          5689 => x"70",
          5690 => x"38",
          5691 => x"05",
          5692 => x"70",
          5693 => x"34",
          5694 => x"eb",
          5695 => x"0d",
          5696 => x"0d",
          5697 => x"54",
          5698 => x"72",
          5699 => x"54",
          5700 => x"51",
          5701 => x"84",
          5702 => x"fc",
          5703 => x"77",
          5704 => x"53",
          5705 => x"05",
          5706 => x"70",
          5707 => x"33",
          5708 => x"ff",
          5709 => x"52",
          5710 => x"2e",
          5711 => x"80",
          5712 => x"71",
          5713 => x"0c",
          5714 => x"04",
          5715 => x"74",
          5716 => x"89",
          5717 => x"2e",
          5718 => x"11",
          5719 => x"52",
          5720 => x"70",
          5721 => x"d8",
          5722 => x"0d",
          5723 => x"82",
          5724 => x"04",
          5725 => x"77",
          5726 => x"70",
          5727 => x"33",
          5728 => x"55",
          5729 => x"ff",
          5730 => x"d8",
          5731 => x"72",
          5732 => x"38",
          5733 => x"72",
          5734 => x"b6",
          5735 => x"d8",
          5736 => x"ff",
          5737 => x"80",
          5738 => x"73",
          5739 => x"55",
          5740 => x"d8",
          5741 => x"0d",
          5742 => x"0d",
          5743 => x"0b",
          5744 => x"56",
          5745 => x"2e",
          5746 => x"81",
          5747 => x"08",
          5748 => x"70",
          5749 => x"33",
          5750 => x"e4",
          5751 => x"d8",
          5752 => x"09",
          5753 => x"38",
          5754 => x"08",
          5755 => x"b4",
          5756 => x"a8",
          5757 => x"a0",
          5758 => x"56",
          5759 => x"27",
          5760 => x"16",
          5761 => x"82",
          5762 => x"06",
          5763 => x"54",
          5764 => x"78",
          5765 => x"33",
          5766 => x"3f",
          5767 => x"5a",
          5768 => x"d8",
          5769 => x"0d",
          5770 => x"0d",
          5771 => x"56",
          5772 => x"b4",
          5773 => x"af",
          5774 => x"fe",
          5775 => x"d6",
          5776 => x"82",
          5777 => x"9f",
          5778 => x"74",
          5779 => x"52",
          5780 => x"51",
          5781 => x"82",
          5782 => x"80",
          5783 => x"ff",
          5784 => x"74",
          5785 => x"76",
          5786 => x"0c",
          5787 => x"04",
          5788 => x"7a",
          5789 => x"fe",
          5790 => x"d6",
          5791 => x"82",
          5792 => x"81",
          5793 => x"33",
          5794 => x"2e",
          5795 => x"80",
          5796 => x"17",
          5797 => x"81",
          5798 => x"06",
          5799 => x"84",
          5800 => x"d6",
          5801 => x"b8",
          5802 => x"56",
          5803 => x"82",
          5804 => x"84",
          5805 => x"fb",
          5806 => x"8b",
          5807 => x"52",
          5808 => x"eb",
          5809 => x"85",
          5810 => x"84",
          5811 => x"fb",
          5812 => x"17",
          5813 => x"a0",
          5814 => x"d3",
          5815 => x"08",
          5816 => x"17",
          5817 => x"3f",
          5818 => x"81",
          5819 => x"19",
          5820 => x"53",
          5821 => x"17",
          5822 => x"c4",
          5823 => x"18",
          5824 => x"80",
          5825 => x"33",
          5826 => x"3f",
          5827 => x"08",
          5828 => x"38",
          5829 => x"82",
          5830 => x"8a",
          5831 => x"fb",
          5832 => x"fe",
          5833 => x"08",
          5834 => x"56",
          5835 => x"74",
          5836 => x"38",
          5837 => x"75",
          5838 => x"16",
          5839 => x"53",
          5840 => x"d8",
          5841 => x"0d",
          5842 => x"0d",
          5843 => x"08",
          5844 => x"81",
          5845 => x"df",
          5846 => x"15",
          5847 => x"d7",
          5848 => x"33",
          5849 => x"82",
          5850 => x"38",
          5851 => x"89",
          5852 => x"2e",
          5853 => x"bf",
          5854 => x"2e",
          5855 => x"81",
          5856 => x"81",
          5857 => x"89",
          5858 => x"08",
          5859 => x"52",
          5860 => x"3f",
          5861 => x"08",
          5862 => x"74",
          5863 => x"14",
          5864 => x"81",
          5865 => x"2a",
          5866 => x"05",
          5867 => x"57",
          5868 => x"f5",
          5869 => x"d8",
          5870 => x"38",
          5871 => x"06",
          5872 => x"33",
          5873 => x"78",
          5874 => x"06",
          5875 => x"5c",
          5876 => x"53",
          5877 => x"38",
          5878 => x"06",
          5879 => x"39",
          5880 => x"a8",
          5881 => x"52",
          5882 => x"bd",
          5883 => x"d8",
          5884 => x"38",
          5885 => x"fe",
          5886 => x"b8",
          5887 => x"cf",
          5888 => x"d8",
          5889 => x"ff",
          5890 => x"39",
          5891 => x"a8",
          5892 => x"52",
          5893 => x"91",
          5894 => x"d8",
          5895 => x"76",
          5896 => x"fc",
          5897 => x"b8",
          5898 => x"ba",
          5899 => x"d8",
          5900 => x"06",
          5901 => x"81",
          5902 => x"d6",
          5903 => x"3d",
          5904 => x"3d",
          5905 => x"7e",
          5906 => x"82",
          5907 => x"27",
          5908 => x"76",
          5909 => x"27",
          5910 => x"75",
          5911 => x"79",
          5912 => x"38",
          5913 => x"89",
          5914 => x"2e",
          5915 => x"80",
          5916 => x"2e",
          5917 => x"81",
          5918 => x"81",
          5919 => x"89",
          5920 => x"08",
          5921 => x"52",
          5922 => x"3f",
          5923 => x"08",
          5924 => x"d8",
          5925 => x"38",
          5926 => x"06",
          5927 => x"81",
          5928 => x"06",
          5929 => x"77",
          5930 => x"2e",
          5931 => x"84",
          5932 => x"06",
          5933 => x"06",
          5934 => x"53",
          5935 => x"81",
          5936 => x"34",
          5937 => x"a8",
          5938 => x"52",
          5939 => x"d9",
          5940 => x"d8",
          5941 => x"d6",
          5942 => x"94",
          5943 => x"ff",
          5944 => x"05",
          5945 => x"54",
          5946 => x"38",
          5947 => x"74",
          5948 => x"06",
          5949 => x"07",
          5950 => x"74",
          5951 => x"39",
          5952 => x"a8",
          5953 => x"52",
          5954 => x"9d",
          5955 => x"d8",
          5956 => x"d6",
          5957 => x"d8",
          5958 => x"ff",
          5959 => x"76",
          5960 => x"06",
          5961 => x"05",
          5962 => x"3f",
          5963 => x"87",
          5964 => x"08",
          5965 => x"51",
          5966 => x"82",
          5967 => x"59",
          5968 => x"08",
          5969 => x"f0",
          5970 => x"82",
          5971 => x"06",
          5972 => x"05",
          5973 => x"54",
          5974 => x"3f",
          5975 => x"08",
          5976 => x"74",
          5977 => x"51",
          5978 => x"81",
          5979 => x"34",
          5980 => x"d8",
          5981 => x"0d",
          5982 => x"0d",
          5983 => x"72",
          5984 => x"56",
          5985 => x"27",
          5986 => x"9c",
          5987 => x"9d",
          5988 => x"2e",
          5989 => x"53",
          5990 => x"51",
          5991 => x"82",
          5992 => x"54",
          5993 => x"08",
          5994 => x"93",
          5995 => x"80",
          5996 => x"54",
          5997 => x"82",
          5998 => x"54",
          5999 => x"74",
          6000 => x"fb",
          6001 => x"d6",
          6002 => x"82",
          6003 => x"80",
          6004 => x"38",
          6005 => x"08",
          6006 => x"38",
          6007 => x"08",
          6008 => x"38",
          6009 => x"52",
          6010 => x"d6",
          6011 => x"d8",
          6012 => x"9c",
          6013 => x"11",
          6014 => x"57",
          6015 => x"74",
          6016 => x"81",
          6017 => x"0c",
          6018 => x"81",
          6019 => x"84",
          6020 => x"55",
          6021 => x"ff",
          6022 => x"54",
          6023 => x"d8",
          6024 => x"0d",
          6025 => x"0d",
          6026 => x"08",
          6027 => x"79",
          6028 => x"17",
          6029 => x"80",
          6030 => x"9c",
          6031 => x"26",
          6032 => x"58",
          6033 => x"52",
          6034 => x"fd",
          6035 => x"74",
          6036 => x"08",
          6037 => x"38",
          6038 => x"08",
          6039 => x"d8",
          6040 => x"82",
          6041 => x"17",
          6042 => x"d8",
          6043 => x"c7",
          6044 => x"94",
          6045 => x"56",
          6046 => x"2e",
          6047 => x"77",
          6048 => x"81",
          6049 => x"38",
          6050 => x"9c",
          6051 => x"26",
          6052 => x"56",
          6053 => x"51",
          6054 => x"80",
          6055 => x"d8",
          6056 => x"09",
          6057 => x"38",
          6058 => x"08",
          6059 => x"d8",
          6060 => x"30",
          6061 => x"80",
          6062 => x"07",
          6063 => x"08",
          6064 => x"55",
          6065 => x"ef",
          6066 => x"d8",
          6067 => x"95",
          6068 => x"08",
          6069 => x"27",
          6070 => x"9c",
          6071 => x"89",
          6072 => x"85",
          6073 => x"db",
          6074 => x"81",
          6075 => x"17",
          6076 => x"89",
          6077 => x"75",
          6078 => x"ac",
          6079 => x"7a",
          6080 => x"3f",
          6081 => x"08",
          6082 => x"38",
          6083 => x"d6",
          6084 => x"2e",
          6085 => x"86",
          6086 => x"d8",
          6087 => x"d6",
          6088 => x"70",
          6089 => x"07",
          6090 => x"7c",
          6091 => x"55",
          6092 => x"f8",
          6093 => x"2e",
          6094 => x"ff",
          6095 => x"55",
          6096 => x"ff",
          6097 => x"76",
          6098 => x"3f",
          6099 => x"08",
          6100 => x"08",
          6101 => x"d6",
          6102 => x"80",
          6103 => x"55",
          6104 => x"94",
          6105 => x"2e",
          6106 => x"53",
          6107 => x"51",
          6108 => x"82",
          6109 => x"55",
          6110 => x"75",
          6111 => x"9c",
          6112 => x"05",
          6113 => x"56",
          6114 => x"26",
          6115 => x"15",
          6116 => x"84",
          6117 => x"07",
          6118 => x"18",
          6119 => x"ff",
          6120 => x"2e",
          6121 => x"39",
          6122 => x"39",
          6123 => x"08",
          6124 => x"81",
          6125 => x"74",
          6126 => x"0c",
          6127 => x"04",
          6128 => x"7a",
          6129 => x"f3",
          6130 => x"d6",
          6131 => x"81",
          6132 => x"d8",
          6133 => x"38",
          6134 => x"51",
          6135 => x"82",
          6136 => x"82",
          6137 => x"b4",
          6138 => x"84",
          6139 => x"52",
          6140 => x"52",
          6141 => x"3f",
          6142 => x"39",
          6143 => x"8a",
          6144 => x"75",
          6145 => x"38",
          6146 => x"19",
          6147 => x"81",
          6148 => x"ed",
          6149 => x"d6",
          6150 => x"2e",
          6151 => x"15",
          6152 => x"70",
          6153 => x"07",
          6154 => x"53",
          6155 => x"75",
          6156 => x"0c",
          6157 => x"04",
          6158 => x"7a",
          6159 => x"58",
          6160 => x"f0",
          6161 => x"80",
          6162 => x"9f",
          6163 => x"80",
          6164 => x"90",
          6165 => x"17",
          6166 => x"aa",
          6167 => x"53",
          6168 => x"88",
          6169 => x"08",
          6170 => x"38",
          6171 => x"53",
          6172 => x"17",
          6173 => x"72",
          6174 => x"fe",
          6175 => x"08",
          6176 => x"80",
          6177 => x"16",
          6178 => x"2b",
          6179 => x"75",
          6180 => x"73",
          6181 => x"f5",
          6182 => x"d6",
          6183 => x"82",
          6184 => x"ff",
          6185 => x"81",
          6186 => x"d8",
          6187 => x"38",
          6188 => x"82",
          6189 => x"26",
          6190 => x"58",
          6191 => x"73",
          6192 => x"39",
          6193 => x"51",
          6194 => x"82",
          6195 => x"98",
          6196 => x"94",
          6197 => x"17",
          6198 => x"58",
          6199 => x"9a",
          6200 => x"81",
          6201 => x"74",
          6202 => x"98",
          6203 => x"83",
          6204 => x"b8",
          6205 => x"0c",
          6206 => x"82",
          6207 => x"8a",
          6208 => x"f8",
          6209 => x"70",
          6210 => x"08",
          6211 => x"57",
          6212 => x"0a",
          6213 => x"38",
          6214 => x"15",
          6215 => x"08",
          6216 => x"72",
          6217 => x"cb",
          6218 => x"ff",
          6219 => x"81",
          6220 => x"13",
          6221 => x"94",
          6222 => x"74",
          6223 => x"85",
          6224 => x"22",
          6225 => x"73",
          6226 => x"38",
          6227 => x"8a",
          6228 => x"05",
          6229 => x"06",
          6230 => x"8a",
          6231 => x"73",
          6232 => x"3f",
          6233 => x"08",
          6234 => x"81",
          6235 => x"d8",
          6236 => x"ff",
          6237 => x"82",
          6238 => x"ff",
          6239 => x"38",
          6240 => x"82",
          6241 => x"26",
          6242 => x"7b",
          6243 => x"98",
          6244 => x"55",
          6245 => x"94",
          6246 => x"73",
          6247 => x"3f",
          6248 => x"08",
          6249 => x"82",
          6250 => x"80",
          6251 => x"38",
          6252 => x"d6",
          6253 => x"2e",
          6254 => x"55",
          6255 => x"08",
          6256 => x"38",
          6257 => x"08",
          6258 => x"fb",
          6259 => x"d6",
          6260 => x"38",
          6261 => x"0c",
          6262 => x"51",
          6263 => x"82",
          6264 => x"98",
          6265 => x"90",
          6266 => x"16",
          6267 => x"15",
          6268 => x"74",
          6269 => x"0c",
          6270 => x"04",
          6271 => x"7b",
          6272 => x"5b",
          6273 => x"52",
          6274 => x"ac",
          6275 => x"d8",
          6276 => x"d6",
          6277 => x"ec",
          6278 => x"d8",
          6279 => x"17",
          6280 => x"51",
          6281 => x"82",
          6282 => x"54",
          6283 => x"08",
          6284 => x"82",
          6285 => x"9c",
          6286 => x"33",
          6287 => x"72",
          6288 => x"09",
          6289 => x"38",
          6290 => x"d6",
          6291 => x"72",
          6292 => x"55",
          6293 => x"53",
          6294 => x"8e",
          6295 => x"56",
          6296 => x"09",
          6297 => x"38",
          6298 => x"d6",
          6299 => x"81",
          6300 => x"fd",
          6301 => x"d6",
          6302 => x"82",
          6303 => x"80",
          6304 => x"38",
          6305 => x"09",
          6306 => x"38",
          6307 => x"82",
          6308 => x"8b",
          6309 => x"fd",
          6310 => x"9a",
          6311 => x"eb",
          6312 => x"d6",
          6313 => x"ff",
          6314 => x"70",
          6315 => x"53",
          6316 => x"09",
          6317 => x"38",
          6318 => x"eb",
          6319 => x"d6",
          6320 => x"2b",
          6321 => x"72",
          6322 => x"0c",
          6323 => x"04",
          6324 => x"77",
          6325 => x"ff",
          6326 => x"9a",
          6327 => x"55",
          6328 => x"76",
          6329 => x"53",
          6330 => x"09",
          6331 => x"38",
          6332 => x"52",
          6333 => x"eb",
          6334 => x"3d",
          6335 => x"3d",
          6336 => x"80",
          6337 => x"70",
          6338 => x"81",
          6339 => x"74",
          6340 => x"56",
          6341 => x"70",
          6342 => x"ff",
          6343 => x"51",
          6344 => x"38",
          6345 => x"d8",
          6346 => x"0d",
          6347 => x"0d",
          6348 => x"59",
          6349 => x"5f",
          6350 => x"70",
          6351 => x"19",
          6352 => x"83",
          6353 => x"19",
          6354 => x"51",
          6355 => x"82",
          6356 => x"5b",
          6357 => x"08",
          6358 => x"9c",
          6359 => x"33",
          6360 => x"86",
          6361 => x"82",
          6362 => x"15",
          6363 => x"70",
          6364 => x"58",
          6365 => x"1a",
          6366 => x"d8",
          6367 => x"81",
          6368 => x"81",
          6369 => x"81",
          6370 => x"d8",
          6371 => x"ae",
          6372 => x"06",
          6373 => x"53",
          6374 => x"53",
          6375 => x"82",
          6376 => x"77",
          6377 => x"56",
          6378 => x"09",
          6379 => x"38",
          6380 => x"7f",
          6381 => x"81",
          6382 => x"ef",
          6383 => x"2e",
          6384 => x"81",
          6385 => x"86",
          6386 => x"06",
          6387 => x"80",
          6388 => x"8d",
          6389 => x"81",
          6390 => x"90",
          6391 => x"1d",
          6392 => x"5d",
          6393 => x"09",
          6394 => x"9c",
          6395 => x"33",
          6396 => x"2e",
          6397 => x"81",
          6398 => x"1e",
          6399 => x"52",
          6400 => x"3f",
          6401 => x"08",
          6402 => x"06",
          6403 => x"f8",
          6404 => x"70",
          6405 => x"8d",
          6406 => x"51",
          6407 => x"58",
          6408 => x"d4",
          6409 => x"05",
          6410 => x"3f",
          6411 => x"08",
          6412 => x"06",
          6413 => x"2e",
          6414 => x"81",
          6415 => x"c8",
          6416 => x"1a",
          6417 => x"75",
          6418 => x"14",
          6419 => x"75",
          6420 => x"2e",
          6421 => x"b0",
          6422 => x"57",
          6423 => x"c1",
          6424 => x"70",
          6425 => x"81",
          6426 => x"55",
          6427 => x"8e",
          6428 => x"fe",
          6429 => x"73",
          6430 => x"80",
          6431 => x"1c",
          6432 => x"06",
          6433 => x"39",
          6434 => x"72",
          6435 => x"7b",
          6436 => x"51",
          6437 => x"82",
          6438 => x"81",
          6439 => x"72",
          6440 => x"38",
          6441 => x"1a",
          6442 => x"80",
          6443 => x"f8",
          6444 => x"d6",
          6445 => x"82",
          6446 => x"89",
          6447 => x"08",
          6448 => x"86",
          6449 => x"98",
          6450 => x"82",
          6451 => x"90",
          6452 => x"f2",
          6453 => x"70",
          6454 => x"80",
          6455 => x"f6",
          6456 => x"d6",
          6457 => x"82",
          6458 => x"83",
          6459 => x"ff",
          6460 => x"ff",
          6461 => x"0c",
          6462 => x"52",
          6463 => x"a9",
          6464 => x"d8",
          6465 => x"d6",
          6466 => x"85",
          6467 => x"08",
          6468 => x"57",
          6469 => x"84",
          6470 => x"39",
          6471 => x"bf",
          6472 => x"ff",
          6473 => x"73",
          6474 => x"75",
          6475 => x"82",
          6476 => x"83",
          6477 => x"06",
          6478 => x"8f",
          6479 => x"73",
          6480 => x"74",
          6481 => x"81",
          6482 => x"38",
          6483 => x"70",
          6484 => x"81",
          6485 => x"55",
          6486 => x"38",
          6487 => x"70",
          6488 => x"54",
          6489 => x"92",
          6490 => x"33",
          6491 => x"06",
          6492 => x"08",
          6493 => x"58",
          6494 => x"7c",
          6495 => x"06",
          6496 => x"8d",
          6497 => x"7d",
          6498 => x"81",
          6499 => x"38",
          6500 => x"9a",
          6501 => x"e5",
          6502 => x"d6",
          6503 => x"ff",
          6504 => x"74",
          6505 => x"76",
          6506 => x"06",
          6507 => x"05",
          6508 => x"75",
          6509 => x"c7",
          6510 => x"77",
          6511 => x"8f",
          6512 => x"d8",
          6513 => x"ff",
          6514 => x"80",
          6515 => x"77",
          6516 => x"80",
          6517 => x"51",
          6518 => x"3f",
          6519 => x"08",
          6520 => x"70",
          6521 => x"81",
          6522 => x"80",
          6523 => x"74",
          6524 => x"08",
          6525 => x"06",
          6526 => x"75",
          6527 => x"75",
          6528 => x"2e",
          6529 => x"b3",
          6530 => x"5b",
          6531 => x"ff",
          6532 => x"33",
          6533 => x"70",
          6534 => x"55",
          6535 => x"2e",
          6536 => x"80",
          6537 => x"77",
          6538 => x"22",
          6539 => x"8b",
          6540 => x"70",
          6541 => x"51",
          6542 => x"81",
          6543 => x"5c",
          6544 => x"93",
          6545 => x"f9",
          6546 => x"d6",
          6547 => x"ff",
          6548 => x"7e",
          6549 => x"ab",
          6550 => x"06",
          6551 => x"38",
          6552 => x"19",
          6553 => x"08",
          6554 => x"3f",
          6555 => x"08",
          6556 => x"38",
          6557 => x"ff",
          6558 => x"0c",
          6559 => x"51",
          6560 => x"82",
          6561 => x"58",
          6562 => x"08",
          6563 => x"e8",
          6564 => x"d6",
          6565 => x"3d",
          6566 => x"3d",
          6567 => x"08",
          6568 => x"81",
          6569 => x"5d",
          6570 => x"73",
          6571 => x"73",
          6572 => x"70",
          6573 => x"5d",
          6574 => x"8d",
          6575 => x"70",
          6576 => x"22",
          6577 => x"f0",
          6578 => x"a0",
          6579 => x"92",
          6580 => x"5f",
          6581 => x"3f",
          6582 => x"05",
          6583 => x"54",
          6584 => x"82",
          6585 => x"c0",
          6586 => x"34",
          6587 => x"1c",
          6588 => x"58",
          6589 => x"52",
          6590 => x"e2",
          6591 => x"27",
          6592 => x"7a",
          6593 => x"70",
          6594 => x"06",
          6595 => x"80",
          6596 => x"74",
          6597 => x"06",
          6598 => x"55",
          6599 => x"81",
          6600 => x"07",
          6601 => x"71",
          6602 => x"81",
          6603 => x"56",
          6604 => x"2e",
          6605 => x"84",
          6606 => x"56",
          6607 => x"76",
          6608 => x"38",
          6609 => x"55",
          6610 => x"05",
          6611 => x"57",
          6612 => x"bf",
          6613 => x"74",
          6614 => x"87",
          6615 => x"76",
          6616 => x"ff",
          6617 => x"2a",
          6618 => x"74",
          6619 => x"3d",
          6620 => x"54",
          6621 => x"34",
          6622 => x"b5",
          6623 => x"54",
          6624 => x"ad",
          6625 => x"70",
          6626 => x"e3",
          6627 => x"d6",
          6628 => x"2e",
          6629 => x"17",
          6630 => x"2e",
          6631 => x"15",
          6632 => x"55",
          6633 => x"89",
          6634 => x"70",
          6635 => x"d0",
          6636 => x"77",
          6637 => x"54",
          6638 => x"16",
          6639 => x"56",
          6640 => x"8a",
          6641 => x"81",
          6642 => x"58",
          6643 => x"78",
          6644 => x"27",
          6645 => x"51",
          6646 => x"82",
          6647 => x"8b",
          6648 => x"5b",
          6649 => x"27",
          6650 => x"87",
          6651 => x"e4",
          6652 => x"38",
          6653 => x"08",
          6654 => x"d8",
          6655 => x"09",
          6656 => x"df",
          6657 => x"cb",
          6658 => x"1b",
          6659 => x"cb",
          6660 => x"81",
          6661 => x"06",
          6662 => x"81",
          6663 => x"2e",
          6664 => x"52",
          6665 => x"fe",
          6666 => x"82",
          6667 => x"19",
          6668 => x"79",
          6669 => x"3f",
          6670 => x"08",
          6671 => x"d8",
          6672 => x"38",
          6673 => x"78",
          6674 => x"d4",
          6675 => x"2b",
          6676 => x"71",
          6677 => x"79",
          6678 => x"3f",
          6679 => x"08",
          6680 => x"d8",
          6681 => x"38",
          6682 => x"f5",
          6683 => x"d6",
          6684 => x"ff",
          6685 => x"1a",
          6686 => x"51",
          6687 => x"82",
          6688 => x"57",
          6689 => x"08",
          6690 => x"8c",
          6691 => x"1b",
          6692 => x"ff",
          6693 => x"5b",
          6694 => x"34",
          6695 => x"17",
          6696 => x"d8",
          6697 => x"34",
          6698 => x"08",
          6699 => x"51",
          6700 => x"77",
          6701 => x"05",
          6702 => x"73",
          6703 => x"2e",
          6704 => x"10",
          6705 => x"81",
          6706 => x"54",
          6707 => x"c7",
          6708 => x"76",
          6709 => x"b9",
          6710 => x"38",
          6711 => x"54",
          6712 => x"8c",
          6713 => x"38",
          6714 => x"ff",
          6715 => x"74",
          6716 => x"22",
          6717 => x"86",
          6718 => x"c0",
          6719 => x"76",
          6720 => x"83",
          6721 => x"52",
          6722 => x"f7",
          6723 => x"d8",
          6724 => x"d6",
          6725 => x"c9",
          6726 => x"59",
          6727 => x"38",
          6728 => x"52",
          6729 => x"81",
          6730 => x"d8",
          6731 => x"d6",
          6732 => x"38",
          6733 => x"d6",
          6734 => x"9c",
          6735 => x"df",
          6736 => x"53",
          6737 => x"9c",
          6738 => x"df",
          6739 => x"1a",
          6740 => x"33",
          6741 => x"55",
          6742 => x"34",
          6743 => x"1d",
          6744 => x"74",
          6745 => x"0c",
          6746 => x"04",
          6747 => x"78",
          6748 => x"12",
          6749 => x"08",
          6750 => x"55",
          6751 => x"94",
          6752 => x"74",
          6753 => x"3f",
          6754 => x"08",
          6755 => x"d8",
          6756 => x"38",
          6757 => x"52",
          6758 => x"8d",
          6759 => x"d8",
          6760 => x"d6",
          6761 => x"38",
          6762 => x"53",
          6763 => x"81",
          6764 => x"34",
          6765 => x"77",
          6766 => x"82",
          6767 => x"52",
          6768 => x"bf",
          6769 => x"d8",
          6770 => x"d6",
          6771 => x"2e",
          6772 => x"84",
          6773 => x"06",
          6774 => x"54",
          6775 => x"d8",
          6776 => x"0d",
          6777 => x"0d",
          6778 => x"08",
          6779 => x"80",
          6780 => x"34",
          6781 => x"80",
          6782 => x"38",
          6783 => x"ff",
          6784 => x"38",
          6785 => x"7f",
          6786 => x"70",
          6787 => x"5b",
          6788 => x"77",
          6789 => x"38",
          6790 => x"70",
          6791 => x"5b",
          6792 => x"97",
          6793 => x"80",
          6794 => x"ff",
          6795 => x"53",
          6796 => x"26",
          6797 => x"5b",
          6798 => x"76",
          6799 => x"81",
          6800 => x"58",
          6801 => x"b5",
          6802 => x"2b",
          6803 => x"80",
          6804 => x"82",
          6805 => x"83",
          6806 => x"55",
          6807 => x"27",
          6808 => x"76",
          6809 => x"74",
          6810 => x"72",
          6811 => x"97",
          6812 => x"55",
          6813 => x"30",
          6814 => x"78",
          6815 => x"72",
          6816 => x"52",
          6817 => x"80",
          6818 => x"80",
          6819 => x"74",
          6820 => x"55",
          6821 => x"80",
          6822 => x"08",
          6823 => x"70",
          6824 => x"54",
          6825 => x"38",
          6826 => x"80",
          6827 => x"79",
          6828 => x"53",
          6829 => x"05",
          6830 => x"82",
          6831 => x"70",
          6832 => x"5a",
          6833 => x"08",
          6834 => x"81",
          6835 => x"53",
          6836 => x"b7",
          6837 => x"2e",
          6838 => x"84",
          6839 => x"55",
          6840 => x"70",
          6841 => x"07",
          6842 => x"54",
          6843 => x"26",
          6844 => x"80",
          6845 => x"ae",
          6846 => x"05",
          6847 => x"17",
          6848 => x"70",
          6849 => x"34",
          6850 => x"8a",
          6851 => x"b5",
          6852 => x"88",
          6853 => x"0b",
          6854 => x"96",
          6855 => x"72",
          6856 => x"76",
          6857 => x"0b",
          6858 => x"81",
          6859 => x"39",
          6860 => x"1a",
          6861 => x"57",
          6862 => x"80",
          6863 => x"18",
          6864 => x"56",
          6865 => x"bf",
          6866 => x"72",
          6867 => x"38",
          6868 => x"8c",
          6869 => x"53",
          6870 => x"87",
          6871 => x"2a",
          6872 => x"72",
          6873 => x"72",
          6874 => x"72",
          6875 => x"38",
          6876 => x"83",
          6877 => x"56",
          6878 => x"70",
          6879 => x"34",
          6880 => x"15",
          6881 => x"33",
          6882 => x"59",
          6883 => x"38",
          6884 => x"05",
          6885 => x"82",
          6886 => x"1c",
          6887 => x"33",
          6888 => x"85",
          6889 => x"19",
          6890 => x"08",
          6891 => x"33",
          6892 => x"9c",
          6893 => x"11",
          6894 => x"aa",
          6895 => x"d8",
          6896 => x"96",
          6897 => x"87",
          6898 => x"d8",
          6899 => x"23",
          6900 => x"d8",
          6901 => x"d6",
          6902 => x"19",
          6903 => x"0d",
          6904 => x"0d",
          6905 => x"41",
          6906 => x"70",
          6907 => x"55",
          6908 => x"83",
          6909 => x"73",
          6910 => x"92",
          6911 => x"2e",
          6912 => x"98",
          6913 => x"1f",
          6914 => x"81",
          6915 => x"64",
          6916 => x"56",
          6917 => x"2e",
          6918 => x"83",
          6919 => x"73",
          6920 => x"70",
          6921 => x"25",
          6922 => x"51",
          6923 => x"38",
          6924 => x"0c",
          6925 => x"51",
          6926 => x"26",
          6927 => x"80",
          6928 => x"34",
          6929 => x"51",
          6930 => x"82",
          6931 => x"56",
          6932 => x"63",
          6933 => x"8c",
          6934 => x"54",
          6935 => x"3d",
          6936 => x"da",
          6937 => x"d6",
          6938 => x"2e",
          6939 => x"83",
          6940 => x"82",
          6941 => x"27",
          6942 => x"10",
          6943 => x"d8",
          6944 => x"55",
          6945 => x"23",
          6946 => x"82",
          6947 => x"83",
          6948 => x"70",
          6949 => x"30",
          6950 => x"71",
          6951 => x"51",
          6952 => x"73",
          6953 => x"80",
          6954 => x"38",
          6955 => x"26",
          6956 => x"52",
          6957 => x"51",
          6958 => x"82",
          6959 => x"81",
          6960 => x"81",
          6961 => x"d7",
          6962 => x"1a",
          6963 => x"23",
          6964 => x"ff",
          6965 => x"15",
          6966 => x"70",
          6967 => x"57",
          6968 => x"09",
          6969 => x"38",
          6970 => x"80",
          6971 => x"30",
          6972 => x"79",
          6973 => x"54",
          6974 => x"74",
          6975 => x"27",
          6976 => x"78",
          6977 => x"81",
          6978 => x"79",
          6979 => x"ae",
          6980 => x"80",
          6981 => x"82",
          6982 => x"06",
          6983 => x"82",
          6984 => x"73",
          6985 => x"81",
          6986 => x"38",
          6987 => x"73",
          6988 => x"81",
          6989 => x"78",
          6990 => x"80",
          6991 => x"0b",
          6992 => x"58",
          6993 => x"78",
          6994 => x"a0",
          6995 => x"70",
          6996 => x"34",
          6997 => x"8a",
          6998 => x"38",
          6999 => x"54",
          7000 => x"34",
          7001 => x"78",
          7002 => x"38",
          7003 => x"fe",
          7004 => x"22",
          7005 => x"72",
          7006 => x"30",
          7007 => x"51",
          7008 => x"56",
          7009 => x"2e",
          7010 => x"87",
          7011 => x"59",
          7012 => x"78",
          7013 => x"55",
          7014 => x"23",
          7015 => x"86",
          7016 => x"39",
          7017 => x"57",
          7018 => x"80",
          7019 => x"83",
          7020 => x"56",
          7021 => x"a0",
          7022 => x"06",
          7023 => x"1d",
          7024 => x"70",
          7025 => x"5d",
          7026 => x"f2",
          7027 => x"38",
          7028 => x"ff",
          7029 => x"ae",
          7030 => x"06",
          7031 => x"83",
          7032 => x"80",
          7033 => x"79",
          7034 => x"70",
          7035 => x"73",
          7036 => x"38",
          7037 => x"fe",
          7038 => x"19",
          7039 => x"2e",
          7040 => x"15",
          7041 => x"55",
          7042 => x"09",
          7043 => x"38",
          7044 => x"52",
          7045 => x"d5",
          7046 => x"70",
          7047 => x"5f",
          7048 => x"70",
          7049 => x"5f",
          7050 => x"80",
          7051 => x"38",
          7052 => x"96",
          7053 => x"32",
          7054 => x"80",
          7055 => x"54",
          7056 => x"8c",
          7057 => x"2e",
          7058 => x"83",
          7059 => x"39",
          7060 => x"5b",
          7061 => x"83",
          7062 => x"7c",
          7063 => x"30",
          7064 => x"80",
          7065 => x"07",
          7066 => x"55",
          7067 => x"a6",
          7068 => x"2e",
          7069 => x"7c",
          7070 => x"38",
          7071 => x"57",
          7072 => x"81",
          7073 => x"5d",
          7074 => x"7c",
          7075 => x"fc",
          7076 => x"ff",
          7077 => x"ff",
          7078 => x"38",
          7079 => x"57",
          7080 => x"75",
          7081 => x"c2",
          7082 => x"d8",
          7083 => x"ff",
          7084 => x"2a",
          7085 => x"51",
          7086 => x"80",
          7087 => x"75",
          7088 => x"82",
          7089 => x"33",
          7090 => x"ff",
          7091 => x"38",
          7092 => x"73",
          7093 => x"38",
          7094 => x"7f",
          7095 => x"c0",
          7096 => x"a0",
          7097 => x"2a",
          7098 => x"75",
          7099 => x"58",
          7100 => x"75",
          7101 => x"38",
          7102 => x"c6",
          7103 => x"cc",
          7104 => x"d8",
          7105 => x"8a",
          7106 => x"77",
          7107 => x"56",
          7108 => x"bf",
          7109 => x"99",
          7110 => x"7b",
          7111 => x"ff",
          7112 => x"73",
          7113 => x"38",
          7114 => x"e0",
          7115 => x"ff",
          7116 => x"55",
          7117 => x"a0",
          7118 => x"74",
          7119 => x"58",
          7120 => x"a0",
          7121 => x"73",
          7122 => x"09",
          7123 => x"38",
          7124 => x"1f",
          7125 => x"2e",
          7126 => x"88",
          7127 => x"2b",
          7128 => x"5c",
          7129 => x"54",
          7130 => x"8d",
          7131 => x"06",
          7132 => x"2e",
          7133 => x"85",
          7134 => x"07",
          7135 => x"2a",
          7136 => x"51",
          7137 => x"38",
          7138 => x"54",
          7139 => x"85",
          7140 => x"07",
          7141 => x"2a",
          7142 => x"51",
          7143 => x"2e",
          7144 => x"88",
          7145 => x"ab",
          7146 => x"51",
          7147 => x"82",
          7148 => x"ab",
          7149 => x"56",
          7150 => x"08",
          7151 => x"38",
          7152 => x"08",
          7153 => x"81",
          7154 => x"38",
          7155 => x"70",
          7156 => x"82",
          7157 => x"54",
          7158 => x"96",
          7159 => x"06",
          7160 => x"2e",
          7161 => x"ff",
          7162 => x"1f",
          7163 => x"80",
          7164 => x"81",
          7165 => x"bb",
          7166 => x"b7",
          7167 => x"2a",
          7168 => x"51",
          7169 => x"38",
          7170 => x"70",
          7171 => x"81",
          7172 => x"55",
          7173 => x"e1",
          7174 => x"08",
          7175 => x"60",
          7176 => x"52",
          7177 => x"ef",
          7178 => x"d8",
          7179 => x"0c",
          7180 => x"75",
          7181 => x"0c",
          7182 => x"04",
          7183 => x"7c",
          7184 => x"08",
          7185 => x"55",
          7186 => x"59",
          7187 => x"81",
          7188 => x"70",
          7189 => x"33",
          7190 => x"52",
          7191 => x"2e",
          7192 => x"ee",
          7193 => x"2e",
          7194 => x"81",
          7195 => x"33",
          7196 => x"81",
          7197 => x"52",
          7198 => x"26",
          7199 => x"14",
          7200 => x"06",
          7201 => x"52",
          7202 => x"80",
          7203 => x"0b",
          7204 => x"59",
          7205 => x"7a",
          7206 => x"70",
          7207 => x"33",
          7208 => x"05",
          7209 => x"9f",
          7210 => x"53",
          7211 => x"89",
          7212 => x"70",
          7213 => x"54",
          7214 => x"12",
          7215 => x"26",
          7216 => x"12",
          7217 => x"06",
          7218 => x"30",
          7219 => x"51",
          7220 => x"2e",
          7221 => x"85",
          7222 => x"be",
          7223 => x"74",
          7224 => x"30",
          7225 => x"9f",
          7226 => x"2a",
          7227 => x"54",
          7228 => x"2e",
          7229 => x"15",
          7230 => x"55",
          7231 => x"ff",
          7232 => x"39",
          7233 => x"86",
          7234 => x"7c",
          7235 => x"51",
          7236 => x"ee",
          7237 => x"70",
          7238 => x"0c",
          7239 => x"04",
          7240 => x"78",
          7241 => x"83",
          7242 => x"0b",
          7243 => x"79",
          7244 => x"d1",
          7245 => x"55",
          7246 => x"08",
          7247 => x"84",
          7248 => x"ce",
          7249 => x"d6",
          7250 => x"ff",
          7251 => x"83",
          7252 => x"d4",
          7253 => x"81",
          7254 => x"38",
          7255 => x"17",
          7256 => x"74",
          7257 => x"09",
          7258 => x"38",
          7259 => x"81",
          7260 => x"30",
          7261 => x"79",
          7262 => x"54",
          7263 => x"74",
          7264 => x"09",
          7265 => x"38",
          7266 => x"c7",
          7267 => x"ee",
          7268 => x"87",
          7269 => x"d8",
          7270 => x"d6",
          7271 => x"2e",
          7272 => x"53",
          7273 => x"52",
          7274 => x"51",
          7275 => x"82",
          7276 => x"55",
          7277 => x"08",
          7278 => x"38",
          7279 => x"82",
          7280 => x"88",
          7281 => x"f2",
          7282 => x"02",
          7283 => x"cb",
          7284 => x"55",
          7285 => x"60",
          7286 => x"3f",
          7287 => x"08",
          7288 => x"80",
          7289 => x"d8",
          7290 => x"84",
          7291 => x"d8",
          7292 => x"82",
          7293 => x"70",
          7294 => x"8c",
          7295 => x"2e",
          7296 => x"73",
          7297 => x"81",
          7298 => x"33",
          7299 => x"80",
          7300 => x"81",
          7301 => x"c6",
          7302 => x"d6",
          7303 => x"ff",
          7304 => x"06",
          7305 => x"98",
          7306 => x"2e",
          7307 => x"74",
          7308 => x"81",
          7309 => x"8a",
          7310 => x"b4",
          7311 => x"39",
          7312 => x"77",
          7313 => x"81",
          7314 => x"33",
          7315 => x"3f",
          7316 => x"08",
          7317 => x"70",
          7318 => x"55",
          7319 => x"86",
          7320 => x"80",
          7321 => x"74",
          7322 => x"81",
          7323 => x"8a",
          7324 => x"fc",
          7325 => x"53",
          7326 => x"fd",
          7327 => x"d6",
          7328 => x"ff",
          7329 => x"82",
          7330 => x"06",
          7331 => x"8c",
          7332 => x"58",
          7333 => x"fa",
          7334 => x"58",
          7335 => x"2e",
          7336 => x"fe",
          7337 => x"be",
          7338 => x"d8",
          7339 => x"78",
          7340 => x"5a",
          7341 => x"90",
          7342 => x"75",
          7343 => x"38",
          7344 => x"3d",
          7345 => x"70",
          7346 => x"08",
          7347 => x"7a",
          7348 => x"38",
          7349 => x"51",
          7350 => x"82",
          7351 => x"81",
          7352 => x"81",
          7353 => x"38",
          7354 => x"83",
          7355 => x"38",
          7356 => x"84",
          7357 => x"38",
          7358 => x"81",
          7359 => x"38",
          7360 => x"51",
          7361 => x"82",
          7362 => x"83",
          7363 => x"53",
          7364 => x"2e",
          7365 => x"84",
          7366 => x"ce",
          7367 => x"af",
          7368 => x"d8",
          7369 => x"ff",
          7370 => x"8d",
          7371 => x"14",
          7372 => x"3f",
          7373 => x"08",
          7374 => x"15",
          7375 => x"14",
          7376 => x"34",
          7377 => x"33",
          7378 => x"81",
          7379 => x"54",
          7380 => x"72",
          7381 => x"98",
          7382 => x"ff",
          7383 => x"29",
          7384 => x"33",
          7385 => x"72",
          7386 => x"72",
          7387 => x"38",
          7388 => x"06",
          7389 => x"2e",
          7390 => x"56",
          7391 => x"80",
          7392 => x"c9",
          7393 => x"d6",
          7394 => x"82",
          7395 => x"88",
          7396 => x"8f",
          7397 => x"56",
          7398 => x"38",
          7399 => x"51",
          7400 => x"82",
          7401 => x"83",
          7402 => x"55",
          7403 => x"80",
          7404 => x"c9",
          7405 => x"d6",
          7406 => x"80",
          7407 => x"c9",
          7408 => x"d6",
          7409 => x"ff",
          7410 => x"8d",
          7411 => x"2e",
          7412 => x"88",
          7413 => x"14",
          7414 => x"05",
          7415 => x"75",
          7416 => x"38",
          7417 => x"52",
          7418 => x"51",
          7419 => x"3f",
          7420 => x"08",
          7421 => x"d8",
          7422 => x"82",
          7423 => x"d6",
          7424 => x"ff",
          7425 => x"26",
          7426 => x"57",
          7427 => x"f5",
          7428 => x"82",
          7429 => x"f5",
          7430 => x"81",
          7431 => x"8d",
          7432 => x"2e",
          7433 => x"82",
          7434 => x"16",
          7435 => x"16",
          7436 => x"70",
          7437 => x"7a",
          7438 => x"0c",
          7439 => x"83",
          7440 => x"06",
          7441 => x"e2",
          7442 => x"83",
          7443 => x"d8",
          7444 => x"ff",
          7445 => x"56",
          7446 => x"38",
          7447 => x"38",
          7448 => x"51",
          7449 => x"82",
          7450 => x"ac",
          7451 => x"82",
          7452 => x"39",
          7453 => x"80",
          7454 => x"38",
          7455 => x"15",
          7456 => x"53",
          7457 => x"8d",
          7458 => x"15",
          7459 => x"76",
          7460 => x"51",
          7461 => x"13",
          7462 => x"8d",
          7463 => x"15",
          7464 => x"cc",
          7465 => x"94",
          7466 => x"0b",
          7467 => x"ff",
          7468 => x"15",
          7469 => x"2e",
          7470 => x"81",
          7471 => x"e8",
          7472 => x"8b",
          7473 => x"d8",
          7474 => x"ff",
          7475 => x"81",
          7476 => x"06",
          7477 => x"81",
          7478 => x"51",
          7479 => x"82",
          7480 => x"80",
          7481 => x"d6",
          7482 => x"15",
          7483 => x"14",
          7484 => x"3f",
          7485 => x"08",
          7486 => x"06",
          7487 => x"d4",
          7488 => x"81",
          7489 => x"38",
          7490 => x"c6",
          7491 => x"d6",
          7492 => x"8b",
          7493 => x"2e",
          7494 => x"b3",
          7495 => x"14",
          7496 => x"3f",
          7497 => x"08",
          7498 => x"e4",
          7499 => x"81",
          7500 => x"84",
          7501 => x"c6",
          7502 => x"d6",
          7503 => x"15",
          7504 => x"14",
          7505 => x"3f",
          7506 => x"08",
          7507 => x"76",
          7508 => x"ee",
          7509 => x"05",
          7510 => x"ee",
          7511 => x"86",
          7512 => x"ee",
          7513 => x"15",
          7514 => x"98",
          7515 => x"56",
          7516 => x"d8",
          7517 => x"0d",
          7518 => x"0d",
          7519 => x"55",
          7520 => x"ba",
          7521 => x"53",
          7522 => x"b2",
          7523 => x"52",
          7524 => x"aa",
          7525 => x"22",
          7526 => x"57",
          7527 => x"2e",
          7528 => x"9a",
          7529 => x"33",
          7530 => x"8d",
          7531 => x"d8",
          7532 => x"52",
          7533 => x"71",
          7534 => x"55",
          7535 => x"53",
          7536 => x"0c",
          7537 => x"d6",
          7538 => x"3d",
          7539 => x"3d",
          7540 => x"05",
          7541 => x"89",
          7542 => x"52",
          7543 => x"3f",
          7544 => x"0b",
          7545 => x"08",
          7546 => x"82",
          7547 => x"84",
          7548 => x"a0",
          7549 => x"55",
          7550 => x"2e",
          7551 => x"74",
          7552 => x"73",
          7553 => x"38",
          7554 => x"78",
          7555 => x"54",
          7556 => x"92",
          7557 => x"89",
          7558 => x"84",
          7559 => x"a7",
          7560 => x"d8",
          7561 => x"82",
          7562 => x"88",
          7563 => x"ea",
          7564 => x"02",
          7565 => x"eb",
          7566 => x"59",
          7567 => x"80",
          7568 => x"38",
          7569 => x"70",
          7570 => x"cc",
          7571 => x"3d",
          7572 => x"58",
          7573 => x"82",
          7574 => x"55",
          7575 => x"08",
          7576 => x"7a",
          7577 => x"8c",
          7578 => x"56",
          7579 => x"82",
          7580 => x"55",
          7581 => x"08",
          7582 => x"80",
          7583 => x"70",
          7584 => x"57",
          7585 => x"83",
          7586 => x"77",
          7587 => x"73",
          7588 => x"ab",
          7589 => x"2e",
          7590 => x"84",
          7591 => x"06",
          7592 => x"51",
          7593 => x"82",
          7594 => x"55",
          7595 => x"b2",
          7596 => x"06",
          7597 => x"b8",
          7598 => x"2a",
          7599 => x"51",
          7600 => x"2e",
          7601 => x"55",
          7602 => x"77",
          7603 => x"74",
          7604 => x"77",
          7605 => x"81",
          7606 => x"73",
          7607 => x"af",
          7608 => x"7a",
          7609 => x"3f",
          7610 => x"08",
          7611 => x"b2",
          7612 => x"8e",
          7613 => x"b7",
          7614 => x"a0",
          7615 => x"34",
          7616 => x"52",
          7617 => x"c8",
          7618 => x"62",
          7619 => x"c3",
          7620 => x"54",
          7621 => x"15",
          7622 => x"2e",
          7623 => x"7a",
          7624 => x"51",
          7625 => x"75",
          7626 => x"d0",
          7627 => x"c9",
          7628 => x"d8",
          7629 => x"d6",
          7630 => x"ca",
          7631 => x"74",
          7632 => x"02",
          7633 => x"70",
          7634 => x"81",
          7635 => x"56",
          7636 => x"86",
          7637 => x"82",
          7638 => x"81",
          7639 => x"06",
          7640 => x"80",
          7641 => x"75",
          7642 => x"73",
          7643 => x"38",
          7644 => x"92",
          7645 => x"7a",
          7646 => x"3f",
          7647 => x"08",
          7648 => x"90",
          7649 => x"55",
          7650 => x"08",
          7651 => x"77",
          7652 => x"81",
          7653 => x"73",
          7654 => x"38",
          7655 => x"07",
          7656 => x"11",
          7657 => x"0c",
          7658 => x"0c",
          7659 => x"52",
          7660 => x"3f",
          7661 => x"08",
          7662 => x"08",
          7663 => x"63",
          7664 => x"5a",
          7665 => x"82",
          7666 => x"82",
          7667 => x"8c",
          7668 => x"7a",
          7669 => x"17",
          7670 => x"23",
          7671 => x"34",
          7672 => x"1a",
          7673 => x"9c",
          7674 => x"0b",
          7675 => x"77",
          7676 => x"81",
          7677 => x"73",
          7678 => x"8d",
          7679 => x"d8",
          7680 => x"81",
          7681 => x"d6",
          7682 => x"1a",
          7683 => x"22",
          7684 => x"7b",
          7685 => x"a8",
          7686 => x"78",
          7687 => x"3f",
          7688 => x"08",
          7689 => x"d8",
          7690 => x"83",
          7691 => x"82",
          7692 => x"ff",
          7693 => x"06",
          7694 => x"55",
          7695 => x"56",
          7696 => x"76",
          7697 => x"51",
          7698 => x"27",
          7699 => x"70",
          7700 => x"5a",
          7701 => x"76",
          7702 => x"74",
          7703 => x"83",
          7704 => x"73",
          7705 => x"38",
          7706 => x"51",
          7707 => x"82",
          7708 => x"85",
          7709 => x"8e",
          7710 => x"2a",
          7711 => x"08",
          7712 => x"0c",
          7713 => x"79",
          7714 => x"73",
          7715 => x"0c",
          7716 => x"04",
          7717 => x"60",
          7718 => x"40",
          7719 => x"80",
          7720 => x"3d",
          7721 => x"78",
          7722 => x"3f",
          7723 => x"08",
          7724 => x"d8",
          7725 => x"91",
          7726 => x"74",
          7727 => x"38",
          7728 => x"c7",
          7729 => x"33",
          7730 => x"87",
          7731 => x"2e",
          7732 => x"95",
          7733 => x"91",
          7734 => x"56",
          7735 => x"81",
          7736 => x"34",
          7737 => x"a3",
          7738 => x"08",
          7739 => x"31",
          7740 => x"27",
          7741 => x"5c",
          7742 => x"82",
          7743 => x"19",
          7744 => x"ff",
          7745 => x"74",
          7746 => x"7e",
          7747 => x"ff",
          7748 => x"2a",
          7749 => x"79",
          7750 => x"87",
          7751 => x"08",
          7752 => x"98",
          7753 => x"78",
          7754 => x"3f",
          7755 => x"08",
          7756 => x"27",
          7757 => x"74",
          7758 => x"a3",
          7759 => x"1a",
          7760 => x"08",
          7761 => x"c3",
          7762 => x"d6",
          7763 => x"2e",
          7764 => x"82",
          7765 => x"1a",
          7766 => x"59",
          7767 => x"2e",
          7768 => x"77",
          7769 => x"11",
          7770 => x"55",
          7771 => x"85",
          7772 => x"31",
          7773 => x"76",
          7774 => x"81",
          7775 => x"ff",
          7776 => x"82",
          7777 => x"fe",
          7778 => x"83",
          7779 => x"56",
          7780 => x"a0",
          7781 => x"08",
          7782 => x"74",
          7783 => x"38",
          7784 => x"b8",
          7785 => x"16",
          7786 => x"89",
          7787 => x"51",
          7788 => x"3f",
          7789 => x"56",
          7790 => x"9c",
          7791 => x"19",
          7792 => x"06",
          7793 => x"31",
          7794 => x"76",
          7795 => x"7b",
          7796 => x"08",
          7797 => x"c0",
          7798 => x"d6",
          7799 => x"ff",
          7800 => x"94",
          7801 => x"ff",
          7802 => x"05",
          7803 => x"ff",
          7804 => x"7b",
          7805 => x"08",
          7806 => x"76",
          7807 => x"08",
          7808 => x"0c",
          7809 => x"f0",
          7810 => x"75",
          7811 => x"0c",
          7812 => x"04",
          7813 => x"60",
          7814 => x"40",
          7815 => x"80",
          7816 => x"3d",
          7817 => x"77",
          7818 => x"3f",
          7819 => x"08",
          7820 => x"d8",
          7821 => x"91",
          7822 => x"74",
          7823 => x"38",
          7824 => x"be",
          7825 => x"33",
          7826 => x"70",
          7827 => x"56",
          7828 => x"74",
          7829 => x"aa",
          7830 => x"82",
          7831 => x"34",
          7832 => x"9e",
          7833 => x"91",
          7834 => x"56",
          7835 => x"94",
          7836 => x"11",
          7837 => x"76",
          7838 => x"75",
          7839 => x"80",
          7840 => x"38",
          7841 => x"70",
          7842 => x"56",
          7843 => x"81",
          7844 => x"11",
          7845 => x"77",
          7846 => x"5c",
          7847 => x"38",
          7848 => x"88",
          7849 => x"74",
          7850 => x"52",
          7851 => x"18",
          7852 => x"51",
          7853 => x"82",
          7854 => x"55",
          7855 => x"08",
          7856 => x"b1",
          7857 => x"2e",
          7858 => x"74",
          7859 => x"95",
          7860 => x"19",
          7861 => x"08",
          7862 => x"88",
          7863 => x"55",
          7864 => x"9c",
          7865 => x"09",
          7866 => x"38",
          7867 => x"bd",
          7868 => x"d6",
          7869 => x"ed",
          7870 => x"08",
          7871 => x"c0",
          7872 => x"d6",
          7873 => x"2e",
          7874 => x"82",
          7875 => x"1b",
          7876 => x"5a",
          7877 => x"2e",
          7878 => x"78",
          7879 => x"11",
          7880 => x"55",
          7881 => x"85",
          7882 => x"31",
          7883 => x"76",
          7884 => x"81",
          7885 => x"ff",
          7886 => x"82",
          7887 => x"fe",
          7888 => x"b4",
          7889 => x"31",
          7890 => x"79",
          7891 => x"84",
          7892 => x"16",
          7893 => x"89",
          7894 => x"52",
          7895 => x"ff",
          7896 => x"7e",
          7897 => x"83",
          7898 => x"89",
          7899 => x"de",
          7900 => x"08",
          7901 => x"26",
          7902 => x"51",
          7903 => x"3f",
          7904 => x"08",
          7905 => x"7e",
          7906 => x"0c",
          7907 => x"19",
          7908 => x"08",
          7909 => x"84",
          7910 => x"57",
          7911 => x"27",
          7912 => x"56",
          7913 => x"52",
          7914 => x"bc",
          7915 => x"d6",
          7916 => x"b1",
          7917 => x"7c",
          7918 => x"08",
          7919 => x"1f",
          7920 => x"ff",
          7921 => x"7e",
          7922 => x"83",
          7923 => x"76",
          7924 => x"17",
          7925 => x"1e",
          7926 => x"18",
          7927 => x"0c",
          7928 => x"58",
          7929 => x"74",
          7930 => x"38",
          7931 => x"8c",
          7932 => x"8a",
          7933 => x"33",
          7934 => x"55",
          7935 => x"34",
          7936 => x"82",
          7937 => x"90",
          7938 => x"f8",
          7939 => x"8b",
          7940 => x"53",
          7941 => x"f2",
          7942 => x"d6",
          7943 => x"82",
          7944 => x"81",
          7945 => x"16",
          7946 => x"2a",
          7947 => x"51",
          7948 => x"80",
          7949 => x"38",
          7950 => x"52",
          7951 => x"bb",
          7952 => x"d6",
          7953 => x"82",
          7954 => x"80",
          7955 => x"16",
          7956 => x"33",
          7957 => x"55",
          7958 => x"34",
          7959 => x"53",
          7960 => x"08",
          7961 => x"3f",
          7962 => x"52",
          7963 => x"ff",
          7964 => x"82",
          7965 => x"52",
          7966 => x"ff",
          7967 => x"76",
          7968 => x"51",
          7969 => x"3f",
          7970 => x"0b",
          7971 => x"78",
          7972 => x"dc",
          7973 => x"d8",
          7974 => x"33",
          7975 => x"55",
          7976 => x"17",
          7977 => x"d6",
          7978 => x"3d",
          7979 => x"3d",
          7980 => x"52",
          7981 => x"3f",
          7982 => x"08",
          7983 => x"d8",
          7984 => x"86",
          7985 => x"52",
          7986 => x"ad",
          7987 => x"d8",
          7988 => x"d6",
          7989 => x"38",
          7990 => x"08",
          7991 => x"82",
          7992 => x"86",
          7993 => x"ff",
          7994 => x"3d",
          7995 => x"3f",
          7996 => x"0b",
          7997 => x"08",
          7998 => x"82",
          7999 => x"82",
          8000 => x"80",
          8001 => x"d6",
          8002 => x"3d",
          8003 => x"3d",
          8004 => x"94",
          8005 => x"52",
          8006 => x"e9",
          8007 => x"d6",
          8008 => x"82",
          8009 => x"80",
          8010 => x"58",
          8011 => x"3d",
          8012 => x"dd",
          8013 => x"d6",
          8014 => x"82",
          8015 => x"bc",
          8016 => x"c7",
          8017 => x"98",
          8018 => x"73",
          8019 => x"38",
          8020 => x"12",
          8021 => x"39",
          8022 => x"33",
          8023 => x"70",
          8024 => x"55",
          8025 => x"2e",
          8026 => x"7f",
          8027 => x"54",
          8028 => x"82",
          8029 => x"98",
          8030 => x"39",
          8031 => x"08",
          8032 => x"81",
          8033 => x"85",
          8034 => x"d6",
          8035 => x"3d",
          8036 => x"a3",
          8037 => x"e1",
          8038 => x"e1",
          8039 => x"5b",
          8040 => x"80",
          8041 => x"3d",
          8042 => x"52",
          8043 => x"51",
          8044 => x"82",
          8045 => x"57",
          8046 => x"08",
          8047 => x"7b",
          8048 => x"0c",
          8049 => x"11",
          8050 => x"3d",
          8051 => x"80",
          8052 => x"54",
          8053 => x"82",
          8054 => x"52",
          8055 => x"70",
          8056 => x"d4",
          8057 => x"d8",
          8058 => x"d6",
          8059 => x"ef",
          8060 => x"3d",
          8061 => x"51",
          8062 => x"3f",
          8063 => x"08",
          8064 => x"d8",
          8065 => x"38",
          8066 => x"08",
          8067 => x"c9",
          8068 => x"d6",
          8069 => x"d6",
          8070 => x"52",
          8071 => x"98",
          8072 => x"d8",
          8073 => x"d6",
          8074 => x"b3",
          8075 => x"74",
          8076 => x"3f",
          8077 => x"08",
          8078 => x"d8",
          8079 => x"80",
          8080 => x"52",
          8081 => x"cf",
          8082 => x"d6",
          8083 => x"a6",
          8084 => x"74",
          8085 => x"3f",
          8086 => x"08",
          8087 => x"d8",
          8088 => x"c9",
          8089 => x"2e",
          8090 => x"86",
          8091 => x"81",
          8092 => x"81",
          8093 => x"df",
          8094 => x"05",
          8095 => x"d6",
          8096 => x"93",
          8097 => x"82",
          8098 => x"56",
          8099 => x"80",
          8100 => x"02",
          8101 => x"55",
          8102 => x"16",
          8103 => x"56",
          8104 => x"38",
          8105 => x"73",
          8106 => x"99",
          8107 => x"2e",
          8108 => x"16",
          8109 => x"ff",
          8110 => x"3d",
          8111 => x"18",
          8112 => x"58",
          8113 => x"33",
          8114 => x"eb",
          8115 => x"80",
          8116 => x"11",
          8117 => x"74",
          8118 => x"39",
          8119 => x"09",
          8120 => x"38",
          8121 => x"e1",
          8122 => x"55",
          8123 => x"34",
          8124 => x"ee",
          8125 => x"84",
          8126 => x"c4",
          8127 => x"70",
          8128 => x"56",
          8129 => x"76",
          8130 => x"81",
          8131 => x"70",
          8132 => x"56",
          8133 => x"82",
          8134 => x"78",
          8135 => x"80",
          8136 => x"27",
          8137 => x"19",
          8138 => x"7a",
          8139 => x"5c",
          8140 => x"55",
          8141 => x"7a",
          8142 => x"5c",
          8143 => x"2e",
          8144 => x"85",
          8145 => x"97",
          8146 => x"3d",
          8147 => x"19",
          8148 => x"33",
          8149 => x"05",
          8150 => x"78",
          8151 => x"80",
          8152 => x"82",
          8153 => x"80",
          8154 => x"04",
          8155 => x"7b",
          8156 => x"fc",
          8157 => x"53",
          8158 => x"fd",
          8159 => x"d8",
          8160 => x"d6",
          8161 => x"fe",
          8162 => x"33",
          8163 => x"f6",
          8164 => x"08",
          8165 => x"27",
          8166 => x"15",
          8167 => x"2a",
          8168 => x"51",
          8169 => x"83",
          8170 => x"94",
          8171 => x"80",
          8172 => x"0c",
          8173 => x"2e",
          8174 => x"79",
          8175 => x"70",
          8176 => x"51",
          8177 => x"2e",
          8178 => x"52",
          8179 => x"fe",
          8180 => x"82",
          8181 => x"ff",
          8182 => x"70",
          8183 => x"fe",
          8184 => x"82",
          8185 => x"73",
          8186 => x"76",
          8187 => x"06",
          8188 => x"0c",
          8189 => x"98",
          8190 => x"58",
          8191 => x"39",
          8192 => x"54",
          8193 => x"73",
          8194 => x"ff",
          8195 => x"82",
          8196 => x"54",
          8197 => x"08",
          8198 => x"9d",
          8199 => x"d8",
          8200 => x"81",
          8201 => x"d6",
          8202 => x"16",
          8203 => x"16",
          8204 => x"2e",
          8205 => x"76",
          8206 => x"de",
          8207 => x"31",
          8208 => x"18",
          8209 => x"90",
          8210 => x"81",
          8211 => x"06",
          8212 => x"56",
          8213 => x"9b",
          8214 => x"74",
          8215 => x"c5",
          8216 => x"d8",
          8217 => x"d6",
          8218 => x"38",
          8219 => x"08",
          8220 => x"73",
          8221 => x"ff",
          8222 => x"82",
          8223 => x"54",
          8224 => x"bf",
          8225 => x"27",
          8226 => x"53",
          8227 => x"08",
          8228 => x"73",
          8229 => x"ff",
          8230 => x"15",
          8231 => x"16",
          8232 => x"ff",
          8233 => x"80",
          8234 => x"73",
          8235 => x"ff",
          8236 => x"82",
          8237 => x"94",
          8238 => x"91",
          8239 => x"53",
          8240 => x"81",
          8241 => x"34",
          8242 => x"39",
          8243 => x"82",
          8244 => x"05",
          8245 => x"08",
          8246 => x"08",
          8247 => x"38",
          8248 => x"0c",
          8249 => x"80",
          8250 => x"72",
          8251 => x"73",
          8252 => x"53",
          8253 => x"8c",
          8254 => x"16",
          8255 => x"38",
          8256 => x"0c",
          8257 => x"82",
          8258 => x"8b",
          8259 => x"f9",
          8260 => x"56",
          8261 => x"80",
          8262 => x"38",
          8263 => x"3d",
          8264 => x"8a",
          8265 => x"51",
          8266 => x"82",
          8267 => x"55",
          8268 => x"08",
          8269 => x"77",
          8270 => x"52",
          8271 => x"a1",
          8272 => x"d8",
          8273 => x"d6",
          8274 => x"c4",
          8275 => x"33",
          8276 => x"55",
          8277 => x"24",
          8278 => x"16",
          8279 => x"2a",
          8280 => x"51",
          8281 => x"80",
          8282 => x"9c",
          8283 => x"77",
          8284 => x"3f",
          8285 => x"08",
          8286 => x"77",
          8287 => x"22",
          8288 => x"74",
          8289 => x"ff",
          8290 => x"82",
          8291 => x"55",
          8292 => x"09",
          8293 => x"38",
          8294 => x"39",
          8295 => x"84",
          8296 => x"0c",
          8297 => x"82",
          8298 => x"89",
          8299 => x"fc",
          8300 => x"87",
          8301 => x"53",
          8302 => x"e7",
          8303 => x"d6",
          8304 => x"38",
          8305 => x"08",
          8306 => x"3d",
          8307 => x"3d",
          8308 => x"89",
          8309 => x"54",
          8310 => x"54",
          8311 => x"82",
          8312 => x"53",
          8313 => x"08",
          8314 => x"74",
          8315 => x"d6",
          8316 => x"73",
          8317 => x"c0",
          8318 => x"d8",
          8319 => x"cb",
          8320 => x"d8",
          8321 => x"51",
          8322 => x"82",
          8323 => x"53",
          8324 => x"08",
          8325 => x"81",
          8326 => x"80",
          8327 => x"82",
          8328 => x"a7",
          8329 => x"73",
          8330 => x"3f",
          8331 => x"51",
          8332 => x"3f",
          8333 => x"08",
          8334 => x"30",
          8335 => x"9f",
          8336 => x"d6",
          8337 => x"51",
          8338 => x"72",
          8339 => x"0c",
          8340 => x"04",
          8341 => x"66",
          8342 => x"89",
          8343 => x"97",
          8344 => x"de",
          8345 => x"d6",
          8346 => x"82",
          8347 => x"b2",
          8348 => x"75",
          8349 => x"3f",
          8350 => x"08",
          8351 => x"d8",
          8352 => x"02",
          8353 => x"33",
          8354 => x"55",
          8355 => x"25",
          8356 => x"55",
          8357 => x"80",
          8358 => x"76",
          8359 => x"ce",
          8360 => x"82",
          8361 => x"95",
          8362 => x"f0",
          8363 => x"65",
          8364 => x"53",
          8365 => x"05",
          8366 => x"51",
          8367 => x"82",
          8368 => x"5b",
          8369 => x"08",
          8370 => x"7c",
          8371 => x"08",
          8372 => x"fe",
          8373 => x"08",
          8374 => x"55",
          8375 => x"91",
          8376 => x"0c",
          8377 => x"81",
          8378 => x"39",
          8379 => x"c9",
          8380 => x"d8",
          8381 => x"55",
          8382 => x"2e",
          8383 => x"80",
          8384 => x"75",
          8385 => x"52",
          8386 => x"05",
          8387 => x"b9",
          8388 => x"d8",
          8389 => x"cf",
          8390 => x"d8",
          8391 => x"cc",
          8392 => x"d8",
          8393 => x"82",
          8394 => x"07",
          8395 => x"05",
          8396 => x"53",
          8397 => x"9c",
          8398 => x"26",
          8399 => x"f9",
          8400 => x"08",
          8401 => x"08",
          8402 => x"98",
          8403 => x"81",
          8404 => x"58",
          8405 => x"3f",
          8406 => x"08",
          8407 => x"d8",
          8408 => x"38",
          8409 => x"77",
          8410 => x"5d",
          8411 => x"74",
          8412 => x"81",
          8413 => x"b8",
          8414 => x"a9",
          8415 => x"d6",
          8416 => x"ff",
          8417 => x"30",
          8418 => x"1b",
          8419 => x"5b",
          8420 => x"39",
          8421 => x"ff",
          8422 => x"82",
          8423 => x"f0",
          8424 => x"30",
          8425 => x"1b",
          8426 => x"5b",
          8427 => x"83",
          8428 => x"58",
          8429 => x"92",
          8430 => x"0c",
          8431 => x"12",
          8432 => x"33",
          8433 => x"54",
          8434 => x"34",
          8435 => x"d8",
          8436 => x"0d",
          8437 => x"0d",
          8438 => x"fc",
          8439 => x"52",
          8440 => x"3f",
          8441 => x"08",
          8442 => x"d8",
          8443 => x"38",
          8444 => x"56",
          8445 => x"38",
          8446 => x"70",
          8447 => x"81",
          8448 => x"55",
          8449 => x"80",
          8450 => x"38",
          8451 => x"54",
          8452 => x"08",
          8453 => x"38",
          8454 => x"82",
          8455 => x"53",
          8456 => x"52",
          8457 => x"b2",
          8458 => x"d6",
          8459 => x"88",
          8460 => x"80",
          8461 => x"17",
          8462 => x"51",
          8463 => x"3f",
          8464 => x"08",
          8465 => x"81",
          8466 => x"81",
          8467 => x"d8",
          8468 => x"09",
          8469 => x"38",
          8470 => x"39",
          8471 => x"77",
          8472 => x"d8",
          8473 => x"08",
          8474 => x"98",
          8475 => x"82",
          8476 => x"52",
          8477 => x"b2",
          8478 => x"d6",
          8479 => x"94",
          8480 => x"18",
          8481 => x"33",
          8482 => x"54",
          8483 => x"34",
          8484 => x"85",
          8485 => x"18",
          8486 => x"74",
          8487 => x"0c",
          8488 => x"04",
          8489 => x"82",
          8490 => x"ff",
          8491 => x"a3",
          8492 => x"93",
          8493 => x"d8",
          8494 => x"d6",
          8495 => x"f9",
          8496 => x"a3",
          8497 => x"96",
          8498 => x"58",
          8499 => x"82",
          8500 => x"55",
          8501 => x"08",
          8502 => x"02",
          8503 => x"33",
          8504 => x"70",
          8505 => x"55",
          8506 => x"73",
          8507 => x"75",
          8508 => x"80",
          8509 => x"c1",
          8510 => x"da",
          8511 => x"81",
          8512 => x"87",
          8513 => x"b1",
          8514 => x"78",
          8515 => x"87",
          8516 => x"d8",
          8517 => x"2a",
          8518 => x"51",
          8519 => x"80",
          8520 => x"38",
          8521 => x"d6",
          8522 => x"15",
          8523 => x"89",
          8524 => x"82",
          8525 => x"5c",
          8526 => x"3d",
          8527 => x"ff",
          8528 => x"82",
          8529 => x"55",
          8530 => x"08",
          8531 => x"82",
          8532 => x"52",
          8533 => x"bb",
          8534 => x"d6",
          8535 => x"82",
          8536 => x"86",
          8537 => x"80",
          8538 => x"d6",
          8539 => x"2e",
          8540 => x"d6",
          8541 => x"c1",
          8542 => x"c7",
          8543 => x"d6",
          8544 => x"d6",
          8545 => x"70",
          8546 => x"08",
          8547 => x"51",
          8548 => x"80",
          8549 => x"73",
          8550 => x"38",
          8551 => x"52",
          8552 => x"af",
          8553 => x"d6",
          8554 => x"74",
          8555 => x"51",
          8556 => x"3f",
          8557 => x"08",
          8558 => x"d6",
          8559 => x"3d",
          8560 => x"3d",
          8561 => x"9a",
          8562 => x"05",
          8563 => x"51",
          8564 => x"82",
          8565 => x"54",
          8566 => x"08",
          8567 => x"78",
          8568 => x"8e",
          8569 => x"58",
          8570 => x"82",
          8571 => x"54",
          8572 => x"08",
          8573 => x"54",
          8574 => x"82",
          8575 => x"84",
          8576 => x"06",
          8577 => x"02",
          8578 => x"33",
          8579 => x"81",
          8580 => x"86",
          8581 => x"fd",
          8582 => x"74",
          8583 => x"70",
          8584 => x"b0",
          8585 => x"d6",
          8586 => x"55",
          8587 => x"d8",
          8588 => x"87",
          8589 => x"d8",
          8590 => x"09",
          8591 => x"38",
          8592 => x"d6",
          8593 => x"2e",
          8594 => x"86",
          8595 => x"81",
          8596 => x"81",
          8597 => x"d6",
          8598 => x"78",
          8599 => x"e0",
          8600 => x"d8",
          8601 => x"d6",
          8602 => x"9f",
          8603 => x"a0",
          8604 => x"51",
          8605 => x"3f",
          8606 => x"0b",
          8607 => x"78",
          8608 => x"80",
          8609 => x"82",
          8610 => x"52",
          8611 => x"51",
          8612 => x"3f",
          8613 => x"b8",
          8614 => x"ff",
          8615 => x"a0",
          8616 => x"11",
          8617 => x"05",
          8618 => x"b2",
          8619 => x"ae",
          8620 => x"15",
          8621 => x"78",
          8622 => x"53",
          8623 => x"90",
          8624 => x"81",
          8625 => x"34",
          8626 => x"bf",
          8627 => x"d6",
          8628 => x"82",
          8629 => x"b3",
          8630 => x"b2",
          8631 => x"96",
          8632 => x"a3",
          8633 => x"53",
          8634 => x"51",
          8635 => x"3f",
          8636 => x"0b",
          8637 => x"78",
          8638 => x"83",
          8639 => x"51",
          8640 => x"3f",
          8641 => x"08",
          8642 => x"80",
          8643 => x"76",
          8644 => x"e5",
          8645 => x"d6",
          8646 => x"3d",
          8647 => x"3d",
          8648 => x"84",
          8649 => x"94",
          8650 => x"aa",
          8651 => x"05",
          8652 => x"51",
          8653 => x"82",
          8654 => x"55",
          8655 => x"08",
          8656 => x"78",
          8657 => x"08",
          8658 => x"70",
          8659 => x"91",
          8660 => x"d8",
          8661 => x"d6",
          8662 => x"be",
          8663 => x"9f",
          8664 => x"a0",
          8665 => x"55",
          8666 => x"38",
          8667 => x"3d",
          8668 => x"3d",
          8669 => x"51",
          8670 => x"3f",
          8671 => x"52",
          8672 => x"52",
          8673 => x"d6",
          8674 => x"08",
          8675 => x"c8",
          8676 => x"d6",
          8677 => x"82",
          8678 => x"97",
          8679 => x"3d",
          8680 => x"81",
          8681 => x"65",
          8682 => x"2e",
          8683 => x"55",
          8684 => x"82",
          8685 => x"84",
          8686 => x"06",
          8687 => x"73",
          8688 => x"d6",
          8689 => x"d8",
          8690 => x"d6",
          8691 => x"ca",
          8692 => x"93",
          8693 => x"ff",
          8694 => x"8d",
          8695 => x"a1",
          8696 => x"af",
          8697 => x"17",
          8698 => x"33",
          8699 => x"70",
          8700 => x"55",
          8701 => x"38",
          8702 => x"54",
          8703 => x"34",
          8704 => x"0b",
          8705 => x"8b",
          8706 => x"84",
          8707 => x"06",
          8708 => x"73",
          8709 => x"e7",
          8710 => x"2e",
          8711 => x"75",
          8712 => x"ff",
          8713 => x"82",
          8714 => x"52",
          8715 => x"a5",
          8716 => x"55",
          8717 => x"08",
          8718 => x"de",
          8719 => x"d8",
          8720 => x"51",
          8721 => x"3f",
          8722 => x"08",
          8723 => x"11",
          8724 => x"82",
          8725 => x"80",
          8726 => x"16",
          8727 => x"ae",
          8728 => x"06",
          8729 => x"53",
          8730 => x"51",
          8731 => x"3f",
          8732 => x"0b",
          8733 => x"87",
          8734 => x"d8",
          8735 => x"77",
          8736 => x"3f",
          8737 => x"08",
          8738 => x"d8",
          8739 => x"78",
          8740 => x"dc",
          8741 => x"d8",
          8742 => x"82",
          8743 => x"aa",
          8744 => x"ec",
          8745 => x"80",
          8746 => x"02",
          8747 => x"e3",
          8748 => x"57",
          8749 => x"3d",
          8750 => x"97",
          8751 => x"87",
          8752 => x"d8",
          8753 => x"d6",
          8754 => x"cf",
          8755 => x"66",
          8756 => x"d0",
          8757 => x"89",
          8758 => x"d8",
          8759 => x"d6",
          8760 => x"38",
          8761 => x"05",
          8762 => x"06",
          8763 => x"73",
          8764 => x"a7",
          8765 => x"09",
          8766 => x"71",
          8767 => x"06",
          8768 => x"55",
          8769 => x"15",
          8770 => x"81",
          8771 => x"34",
          8772 => x"a2",
          8773 => x"d6",
          8774 => x"74",
          8775 => x"0c",
          8776 => x"04",
          8777 => x"65",
          8778 => x"94",
          8779 => x"52",
          8780 => x"d1",
          8781 => x"d6",
          8782 => x"82",
          8783 => x"80",
          8784 => x"58",
          8785 => x"3d",
          8786 => x"c5",
          8787 => x"d6",
          8788 => x"82",
          8789 => x"b4",
          8790 => x"c7",
          8791 => x"a0",
          8792 => x"55",
          8793 => x"84",
          8794 => x"17",
          8795 => x"2b",
          8796 => x"96",
          8797 => x"9e",
          8798 => x"54",
          8799 => x"15",
          8800 => x"ff",
          8801 => x"82",
          8802 => x"55",
          8803 => x"d8",
          8804 => x"0d",
          8805 => x"0d",
          8806 => x"5a",
          8807 => x"3d",
          8808 => x"9a",
          8809 => x"9f",
          8810 => x"d8",
          8811 => x"d8",
          8812 => x"82",
          8813 => x"07",
          8814 => x"55",
          8815 => x"2e",
          8816 => x"81",
          8817 => x"55",
          8818 => x"2e",
          8819 => x"7b",
          8820 => x"80",
          8821 => x"70",
          8822 => x"ac",
          8823 => x"d6",
          8824 => x"82",
          8825 => x"80",
          8826 => x"52",
          8827 => x"b2",
          8828 => x"d6",
          8829 => x"82",
          8830 => x"bf",
          8831 => x"d8",
          8832 => x"d8",
          8833 => x"59",
          8834 => x"81",
          8835 => x"56",
          8836 => x"33",
          8837 => x"16",
          8838 => x"27",
          8839 => x"56",
          8840 => x"80",
          8841 => x"80",
          8842 => x"ff",
          8843 => x"70",
          8844 => x"56",
          8845 => x"e8",
          8846 => x"76",
          8847 => x"81",
          8848 => x"80",
          8849 => x"57",
          8850 => x"78",
          8851 => x"51",
          8852 => x"2e",
          8853 => x"73",
          8854 => x"38",
          8855 => x"08",
          8856 => x"9f",
          8857 => x"d6",
          8858 => x"82",
          8859 => x"a7",
          8860 => x"33",
          8861 => x"c3",
          8862 => x"2e",
          8863 => x"e4",
          8864 => x"2e",
          8865 => x"56",
          8866 => x"05",
          8867 => x"d6",
          8868 => x"d8",
          8869 => x"76",
          8870 => x"0c",
          8871 => x"04",
          8872 => x"82",
          8873 => x"ff",
          8874 => x"9d",
          8875 => x"97",
          8876 => x"d8",
          8877 => x"d8",
          8878 => x"82",
          8879 => x"82",
          8880 => x"53",
          8881 => x"3d",
          8882 => x"ff",
          8883 => x"73",
          8884 => x"51",
          8885 => x"74",
          8886 => x"38",
          8887 => x"3d",
          8888 => x"90",
          8889 => x"d8",
          8890 => x"ff",
          8891 => x"38",
          8892 => x"08",
          8893 => x"3f",
          8894 => x"82",
          8895 => x"51",
          8896 => x"82",
          8897 => x"83",
          8898 => x"55",
          8899 => x"a3",
          8900 => x"82",
          8901 => x"ff",
          8902 => x"82",
          8903 => x"93",
          8904 => x"75",
          8905 => x"75",
          8906 => x"38",
          8907 => x"76",
          8908 => x"86",
          8909 => x"39",
          8910 => x"27",
          8911 => x"88",
          8912 => x"77",
          8913 => x"59",
          8914 => x"56",
          8915 => x"81",
          8916 => x"81",
          8917 => x"33",
          8918 => x"73",
          8919 => x"fe",
          8920 => x"33",
          8921 => x"73",
          8922 => x"81",
          8923 => x"80",
          8924 => x"02",
          8925 => x"75",
          8926 => x"51",
          8927 => x"2e",
          8928 => x"87",
          8929 => x"56",
          8930 => x"78",
          8931 => x"80",
          8932 => x"70",
          8933 => x"a9",
          8934 => x"d6",
          8935 => x"82",
          8936 => x"80",
          8937 => x"52",
          8938 => x"af",
          8939 => x"d6",
          8940 => x"82",
          8941 => x"8d",
          8942 => x"c4",
          8943 => x"e5",
          8944 => x"c6",
          8945 => x"d8",
          8946 => x"09",
          8947 => x"cc",
          8948 => x"75",
          8949 => x"c4",
          8950 => x"74",
          8951 => x"9c",
          8952 => x"d8",
          8953 => x"d6",
          8954 => x"38",
          8955 => x"d6",
          8956 => x"66",
          8957 => x"89",
          8958 => x"88",
          8959 => x"34",
          8960 => x"52",
          8961 => x"99",
          8962 => x"54",
          8963 => x"15",
          8964 => x"ff",
          8965 => x"82",
          8966 => x"54",
          8967 => x"82",
          8968 => x"9c",
          8969 => x"f2",
          8970 => x"62",
          8971 => x"80",
          8972 => x"93",
          8973 => x"55",
          8974 => x"5e",
          8975 => x"3f",
          8976 => x"08",
          8977 => x"d8",
          8978 => x"38",
          8979 => x"58",
          8980 => x"38",
          8981 => x"97",
          8982 => x"08",
          8983 => x"38",
          8984 => x"70",
          8985 => x"81",
          8986 => x"55",
          8987 => x"87",
          8988 => x"39",
          8989 => x"90",
          8990 => x"82",
          8991 => x"8a",
          8992 => x"89",
          8993 => x"7f",
          8994 => x"56",
          8995 => x"3f",
          8996 => x"06",
          8997 => x"72",
          8998 => x"82",
          8999 => x"05",
          9000 => x"7c",
          9001 => x"55",
          9002 => x"27",
          9003 => x"16",
          9004 => x"83",
          9005 => x"76",
          9006 => x"80",
          9007 => x"79",
          9008 => x"85",
          9009 => x"7f",
          9010 => x"14",
          9011 => x"83",
          9012 => x"82",
          9013 => x"81",
          9014 => x"38",
          9015 => x"08",
          9016 => x"95",
          9017 => x"d8",
          9018 => x"81",
          9019 => x"7b",
          9020 => x"06",
          9021 => x"39",
          9022 => x"56",
          9023 => x"09",
          9024 => x"b9",
          9025 => x"80",
          9026 => x"80",
          9027 => x"78",
          9028 => x"7a",
          9029 => x"38",
          9030 => x"73",
          9031 => x"81",
          9032 => x"ff",
          9033 => x"74",
          9034 => x"ff",
          9035 => x"82",
          9036 => x"58",
          9037 => x"08",
          9038 => x"74",
          9039 => x"16",
          9040 => x"73",
          9041 => x"39",
          9042 => x"7e",
          9043 => x"0c",
          9044 => x"2e",
          9045 => x"88",
          9046 => x"8c",
          9047 => x"1a",
          9048 => x"07",
          9049 => x"1b",
          9050 => x"08",
          9051 => x"16",
          9052 => x"75",
          9053 => x"38",
          9054 => x"94",
          9055 => x"15",
          9056 => x"54",
          9057 => x"34",
          9058 => x"82",
          9059 => x"90",
          9060 => x"e9",
          9061 => x"6d",
          9062 => x"80",
          9063 => x"9d",
          9064 => x"5c",
          9065 => x"3f",
          9066 => x"0b",
          9067 => x"08",
          9068 => x"38",
          9069 => x"08",
          9070 => x"ee",
          9071 => x"08",
          9072 => x"80",
          9073 => x"80",
          9074 => x"d6",
          9075 => x"ff",
          9076 => x"52",
          9077 => x"8e",
          9078 => x"d6",
          9079 => x"ff",
          9080 => x"06",
          9081 => x"56",
          9082 => x"38",
          9083 => x"70",
          9084 => x"55",
          9085 => x"8b",
          9086 => x"3d",
          9087 => x"83",
          9088 => x"ff",
          9089 => x"82",
          9090 => x"99",
          9091 => x"74",
          9092 => x"38",
          9093 => x"80",
          9094 => x"ff",
          9095 => x"55",
          9096 => x"83",
          9097 => x"78",
          9098 => x"38",
          9099 => x"26",
          9100 => x"81",
          9101 => x"8b",
          9102 => x"79",
          9103 => x"80",
          9104 => x"93",
          9105 => x"39",
          9106 => x"6e",
          9107 => x"89",
          9108 => x"48",
          9109 => x"83",
          9110 => x"61",
          9111 => x"25",
          9112 => x"55",
          9113 => x"8a",
          9114 => x"3d",
          9115 => x"81",
          9116 => x"ff",
          9117 => x"81",
          9118 => x"d8",
          9119 => x"38",
          9120 => x"70",
          9121 => x"d6",
          9122 => x"56",
          9123 => x"38",
          9124 => x"55",
          9125 => x"75",
          9126 => x"38",
          9127 => x"70",
          9128 => x"ff",
          9129 => x"83",
          9130 => x"78",
          9131 => x"89",
          9132 => x"81",
          9133 => x"06",
          9134 => x"80",
          9135 => x"77",
          9136 => x"74",
          9137 => x"8d",
          9138 => x"06",
          9139 => x"2e",
          9140 => x"77",
          9141 => x"93",
          9142 => x"74",
          9143 => x"cb",
          9144 => x"7d",
          9145 => x"81",
          9146 => x"38",
          9147 => x"66",
          9148 => x"81",
          9149 => x"88",
          9150 => x"74",
          9151 => x"38",
          9152 => x"98",
          9153 => x"88",
          9154 => x"82",
          9155 => x"57",
          9156 => x"80",
          9157 => x"76",
          9158 => x"38",
          9159 => x"51",
          9160 => x"3f",
          9161 => x"08",
          9162 => x"87",
          9163 => x"2a",
          9164 => x"5c",
          9165 => x"d6",
          9166 => x"80",
          9167 => x"44",
          9168 => x"0a",
          9169 => x"ec",
          9170 => x"39",
          9171 => x"66",
          9172 => x"81",
          9173 => x"f8",
          9174 => x"74",
          9175 => x"38",
          9176 => x"98",
          9177 => x"f8",
          9178 => x"82",
          9179 => x"57",
          9180 => x"80",
          9181 => x"76",
          9182 => x"38",
          9183 => x"51",
          9184 => x"3f",
          9185 => x"08",
          9186 => x"57",
          9187 => x"08",
          9188 => x"96",
          9189 => x"82",
          9190 => x"10",
          9191 => x"08",
          9192 => x"72",
          9193 => x"59",
          9194 => x"ff",
          9195 => x"5d",
          9196 => x"44",
          9197 => x"11",
          9198 => x"70",
          9199 => x"71",
          9200 => x"06",
          9201 => x"52",
          9202 => x"40",
          9203 => x"09",
          9204 => x"38",
          9205 => x"18",
          9206 => x"39",
          9207 => x"79",
          9208 => x"70",
          9209 => x"58",
          9210 => x"76",
          9211 => x"38",
          9212 => x"7d",
          9213 => x"70",
          9214 => x"55",
          9215 => x"3f",
          9216 => x"08",
          9217 => x"2e",
          9218 => x"9b",
          9219 => x"d8",
          9220 => x"f5",
          9221 => x"38",
          9222 => x"38",
          9223 => x"59",
          9224 => x"38",
          9225 => x"7d",
          9226 => x"81",
          9227 => x"38",
          9228 => x"0b",
          9229 => x"08",
          9230 => x"78",
          9231 => x"1a",
          9232 => x"c0",
          9233 => x"74",
          9234 => x"39",
          9235 => x"55",
          9236 => x"8f",
          9237 => x"fd",
          9238 => x"d6",
          9239 => x"f5",
          9240 => x"78",
          9241 => x"79",
          9242 => x"80",
          9243 => x"f1",
          9244 => x"39",
          9245 => x"81",
          9246 => x"06",
          9247 => x"55",
          9248 => x"27",
          9249 => x"81",
          9250 => x"56",
          9251 => x"38",
          9252 => x"80",
          9253 => x"ff",
          9254 => x"8b",
          9255 => x"90",
          9256 => x"ff",
          9257 => x"84",
          9258 => x"1b",
          9259 => x"e1",
          9260 => x"1c",
          9261 => x"ff",
          9262 => x"8e",
          9263 => x"8f",
          9264 => x"0b",
          9265 => x"7d",
          9266 => x"30",
          9267 => x"84",
          9268 => x"51",
          9269 => x"51",
          9270 => x"3f",
          9271 => x"83",
          9272 => x"90",
          9273 => x"ff",
          9274 => x"93",
          9275 => x"8f",
          9276 => x"39",
          9277 => x"1b",
          9278 => x"b3",
          9279 => x"95",
          9280 => x"52",
          9281 => x"ff",
          9282 => x"81",
          9283 => x"1b",
          9284 => x"fd",
          9285 => x"9c",
          9286 => x"8f",
          9287 => x"83",
          9288 => x"06",
          9289 => x"82",
          9290 => x"52",
          9291 => x"51",
          9292 => x"3f",
          9293 => x"1b",
          9294 => x"f3",
          9295 => x"ac",
          9296 => x"8e",
          9297 => x"52",
          9298 => x"ff",
          9299 => x"86",
          9300 => x"51",
          9301 => x"3f",
          9302 => x"80",
          9303 => x"a9",
          9304 => x"1c",
          9305 => x"82",
          9306 => x"80",
          9307 => x"ae",
          9308 => x"b2",
          9309 => x"1b",
          9310 => x"b3",
          9311 => x"ff",
          9312 => x"96",
          9313 => x"8e",
          9314 => x"80",
          9315 => x"34",
          9316 => x"1c",
          9317 => x"82",
          9318 => x"ab",
          9319 => x"8e",
          9320 => x"d4",
          9321 => x"fe",
          9322 => x"59",
          9323 => x"3f",
          9324 => x"53",
          9325 => x"51",
          9326 => x"3f",
          9327 => x"d6",
          9328 => x"e7",
          9329 => x"2e",
          9330 => x"80",
          9331 => x"54",
          9332 => x"53",
          9333 => x"51",
          9334 => x"3f",
          9335 => x"80",
          9336 => x"ff",
          9337 => x"84",
          9338 => x"d2",
          9339 => x"ff",
          9340 => x"86",
          9341 => x"f2",
          9342 => x"1b",
          9343 => x"af",
          9344 => x"52",
          9345 => x"51",
          9346 => x"3f",
          9347 => x"ec",
          9348 => x"8d",
          9349 => x"d4",
          9350 => x"51",
          9351 => x"3f",
          9352 => x"87",
          9353 => x"52",
          9354 => x"89",
          9355 => x"54",
          9356 => x"7a",
          9357 => x"ff",
          9358 => x"65",
          9359 => x"7a",
          9360 => x"bd",
          9361 => x"80",
          9362 => x"2e",
          9363 => x"9a",
          9364 => x"7a",
          9365 => x"d7",
          9366 => x"84",
          9367 => x"8c",
          9368 => x"0a",
          9369 => x"51",
          9370 => x"ff",
          9371 => x"7d",
          9372 => x"38",
          9373 => x"52",
          9374 => x"8c",
          9375 => x"55",
          9376 => x"62",
          9377 => x"74",
          9378 => x"75",
          9379 => x"7e",
          9380 => x"ac",
          9381 => x"d8",
          9382 => x"38",
          9383 => x"82",
          9384 => x"52",
          9385 => x"8c",
          9386 => x"16",
          9387 => x"56",
          9388 => x"38",
          9389 => x"77",
          9390 => x"8d",
          9391 => x"7d",
          9392 => x"38",
          9393 => x"57",
          9394 => x"83",
          9395 => x"76",
          9396 => x"7a",
          9397 => x"ff",
          9398 => x"82",
          9399 => x"81",
          9400 => x"16",
          9401 => x"56",
          9402 => x"38",
          9403 => x"83",
          9404 => x"86",
          9405 => x"ff",
          9406 => x"38",
          9407 => x"82",
          9408 => x"81",
          9409 => x"06",
          9410 => x"fe",
          9411 => x"53",
          9412 => x"51",
          9413 => x"3f",
          9414 => x"52",
          9415 => x"8a",
          9416 => x"be",
          9417 => x"75",
          9418 => x"81",
          9419 => x"0b",
          9420 => x"77",
          9421 => x"75",
          9422 => x"60",
          9423 => x"80",
          9424 => x"75",
          9425 => x"e8",
          9426 => x"85",
          9427 => x"d6",
          9428 => x"2a",
          9429 => x"75",
          9430 => x"82",
          9431 => x"87",
          9432 => x"52",
          9433 => x"51",
          9434 => x"3f",
          9435 => x"ca",
          9436 => x"8a",
          9437 => x"54",
          9438 => x"52",
          9439 => x"86",
          9440 => x"56",
          9441 => x"08",
          9442 => x"53",
          9443 => x"51",
          9444 => x"3f",
          9445 => x"d6",
          9446 => x"38",
          9447 => x"56",
          9448 => x"56",
          9449 => x"d6",
          9450 => x"75",
          9451 => x"0c",
          9452 => x"04",
          9453 => x"7d",
          9454 => x"80",
          9455 => x"05",
          9456 => x"76",
          9457 => x"38",
          9458 => x"11",
          9459 => x"53",
          9460 => x"79",
          9461 => x"3f",
          9462 => x"09",
          9463 => x"38",
          9464 => x"55",
          9465 => x"db",
          9466 => x"70",
          9467 => x"34",
          9468 => x"74",
          9469 => x"81",
          9470 => x"80",
          9471 => x"55",
          9472 => x"76",
          9473 => x"d6",
          9474 => x"3d",
          9475 => x"3d",
          9476 => x"84",
          9477 => x"33",
          9478 => x"8a",
          9479 => x"06",
          9480 => x"52",
          9481 => x"3f",
          9482 => x"56",
          9483 => x"be",
          9484 => x"08",
          9485 => x"05",
          9486 => x"75",
          9487 => x"56",
          9488 => x"a1",
          9489 => x"fc",
          9490 => x"53",
          9491 => x"76",
          9492 => x"c0",
          9493 => x"32",
          9494 => x"72",
          9495 => x"70",
          9496 => x"56",
          9497 => x"18",
          9498 => x"88",
          9499 => x"3d",
          9500 => x"3d",
          9501 => x"11",
          9502 => x"80",
          9503 => x"38",
          9504 => x"05",
          9505 => x"8c",
          9506 => x"08",
          9507 => x"3f",
          9508 => x"08",
          9509 => x"16",
          9510 => x"09",
          9511 => x"38",
          9512 => x"55",
          9513 => x"55",
          9514 => x"d8",
          9515 => x"0d",
          9516 => x"0d",
          9517 => x"cc",
          9518 => x"73",
          9519 => x"c1",
          9520 => x"0c",
          9521 => x"04",
          9522 => x"02",
          9523 => x"33",
          9524 => x"3d",
          9525 => x"54",
          9526 => x"52",
          9527 => x"ae",
          9528 => x"ff",
          9529 => x"3d",
          9530 => x"3d",
          9531 => x"84",
          9532 => x"22",
          9533 => x"52",
          9534 => x"26",
          9535 => x"83",
          9536 => x"52",
          9537 => x"83",
          9538 => x"27",
          9539 => x"b5",
          9540 => x"06",
          9541 => x"80",
          9542 => x"82",
          9543 => x"51",
          9544 => x"9c",
          9545 => x"70",
          9546 => x"06",
          9547 => x"80",
          9548 => x"38",
          9549 => x"c9",
          9550 => x"22",
          9551 => x"39",
          9552 => x"70",
          9553 => x"53",
          9554 => x"d6",
          9555 => x"3d",
          9556 => x"3d",
          9557 => x"05",
          9558 => x"05",
          9559 => x"53",
          9560 => x"70",
          9561 => x"85",
          9562 => x"9a",
          9563 => x"b5",
          9564 => x"06",
          9565 => x"81",
          9566 => x"38",
          9567 => x"c7",
          9568 => x"22",
          9569 => x"82",
          9570 => x"84",
          9571 => x"fb",
          9572 => x"51",
          9573 => x"ff",
          9574 => x"38",
          9575 => x"ff",
          9576 => x"98",
          9577 => x"ff",
          9578 => x"38",
          9579 => x"56",
          9580 => x"05",
          9581 => x"30",
          9582 => x"72",
          9583 => x"51",
          9584 => x"80",
          9585 => x"70",
          9586 => x"22",
          9587 => x"71",
          9588 => x"70",
          9589 => x"55",
          9590 => x"25",
          9591 => x"73",
          9592 => x"dc",
          9593 => x"29",
          9594 => x"05",
          9595 => x"04",
          9596 => x"10",
          9597 => x"22",
          9598 => x"80",
          9599 => x"75",
          9600 => x"72",
          9601 => x"51",
          9602 => x"12",
          9603 => x"e0",
          9604 => x"39",
          9605 => x"95",
          9606 => x"51",
          9607 => x"12",
          9608 => x"ff",
          9609 => x"85",
          9610 => x"12",
          9611 => x"ff",
          9612 => x"8c",
          9613 => x"f8",
          9614 => x"16",
          9615 => x"39",
          9616 => x"82",
          9617 => x"87",
          9618 => x"00",
          9619 => x"ff",
          9620 => x"00",
          9621 => x"ff",
          9622 => x"ff",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"69",
          9769 => x"00",
          9770 => x"69",
          9771 => x"6c",
          9772 => x"69",
          9773 => x"00",
          9774 => x"6c",
          9775 => x"00",
          9776 => x"65",
          9777 => x"00",
          9778 => x"63",
          9779 => x"72",
          9780 => x"63",
          9781 => x"00",
          9782 => x"64",
          9783 => x"00",
          9784 => x"64",
          9785 => x"00",
          9786 => x"65",
          9787 => x"65",
          9788 => x"65",
          9789 => x"69",
          9790 => x"69",
          9791 => x"66",
          9792 => x"66",
          9793 => x"61",
          9794 => x"00",
          9795 => x"6d",
          9796 => x"65",
          9797 => x"72",
          9798 => x"65",
          9799 => x"00",
          9800 => x"6e",
          9801 => x"00",
          9802 => x"65",
          9803 => x"00",
          9804 => x"62",
          9805 => x"63",
          9806 => x"62",
          9807 => x"63",
          9808 => x"69",
          9809 => x"00",
          9810 => x"64",
          9811 => x"69",
          9812 => x"45",
          9813 => x"72",
          9814 => x"6e",
          9815 => x"6e",
          9816 => x"65",
          9817 => x"72",
          9818 => x"69",
          9819 => x"6e",
          9820 => x"72",
          9821 => x"79",
          9822 => x"6f",
          9823 => x"6c",
          9824 => x"6f",
          9825 => x"2e",
          9826 => x"6f",
          9827 => x"74",
          9828 => x"6f",
          9829 => x"2e",
          9830 => x"6e",
          9831 => x"69",
          9832 => x"69",
          9833 => x"61",
          9834 => x"00",
          9835 => x"63",
          9836 => x"73",
          9837 => x"6e",
          9838 => x"2e",
          9839 => x"69",
          9840 => x"61",
          9841 => x"61",
          9842 => x"65",
          9843 => x"74",
          9844 => x"00",
          9845 => x"69",
          9846 => x"68",
          9847 => x"6c",
          9848 => x"6e",
          9849 => x"69",
          9850 => x"00",
          9851 => x"44",
          9852 => x"20",
          9853 => x"74",
          9854 => x"72",
          9855 => x"63",
          9856 => x"2e",
          9857 => x"72",
          9858 => x"20",
          9859 => x"62",
          9860 => x"69",
          9861 => x"6e",
          9862 => x"69",
          9863 => x"00",
          9864 => x"69",
          9865 => x"6e",
          9866 => x"65",
          9867 => x"6c",
          9868 => x"00",
          9869 => x"6f",
          9870 => x"6d",
          9871 => x"69",
          9872 => x"20",
          9873 => x"65",
          9874 => x"74",
          9875 => x"66",
          9876 => x"64",
          9877 => x"20",
          9878 => x"6b",
          9879 => x"6f",
          9880 => x"74",
          9881 => x"6f",
          9882 => x"64",
          9883 => x"69",
          9884 => x"75",
          9885 => x"6f",
          9886 => x"61",
          9887 => x"6e",
          9888 => x"6e",
          9889 => x"6c",
          9890 => x"00",
          9891 => x"69",
          9892 => x"69",
          9893 => x"6f",
          9894 => x"64",
          9895 => x"6e",
          9896 => x"66",
          9897 => x"65",
          9898 => x"6d",
          9899 => x"72",
          9900 => x"00",
          9901 => x"6f",
          9902 => x"61",
          9903 => x"6f",
          9904 => x"20",
          9905 => x"65",
          9906 => x"00",
          9907 => x"61",
          9908 => x"65",
          9909 => x"73",
          9910 => x"63",
          9911 => x"65",
          9912 => x"00",
          9913 => x"75",
          9914 => x"73",
          9915 => x"00",
          9916 => x"6e",
          9917 => x"77",
          9918 => x"72",
          9919 => x"2e",
          9920 => x"25",
          9921 => x"62",
          9922 => x"73",
          9923 => x"20",
          9924 => x"25",
          9925 => x"62",
          9926 => x"73",
          9927 => x"63",
          9928 => x"00",
          9929 => x"65",
          9930 => x"00",
          9931 => x"3d",
          9932 => x"6c",
          9933 => x"31",
          9934 => x"38",
          9935 => x"20",
          9936 => x"30",
          9937 => x"2c",
          9938 => x"4f",
          9939 => x"30",
          9940 => x"20",
          9941 => x"6c",
          9942 => x"30",
          9943 => x"0a",
          9944 => x"30",
          9945 => x"00",
          9946 => x"20",
          9947 => x"30",
          9948 => x"00",
          9949 => x"20",
          9950 => x"20",
          9951 => x"00",
          9952 => x"30",
          9953 => x"00",
          9954 => x"20",
          9955 => x"7c",
          9956 => x"00",
          9957 => x"4f",
          9958 => x"2a",
          9959 => x"73",
          9960 => x"00",
          9961 => x"35",
          9962 => x"2f",
          9963 => x"30",
          9964 => x"31",
          9965 => x"66",
          9966 => x"5a",
          9967 => x"20",
          9968 => x"20",
          9969 => x"78",
          9970 => x"73",
          9971 => x"20",
          9972 => x"0a",
          9973 => x"50",
          9974 => x"6e",
          9975 => x"72",
          9976 => x"20",
          9977 => x"64",
          9978 => x"00",
          9979 => x"69",
          9980 => x"20",
          9981 => x"65",
          9982 => x"70",
          9983 => x"53",
          9984 => x"6e",
          9985 => x"72",
          9986 => x"00",
          9987 => x"4f",
          9988 => x"20",
          9989 => x"69",
          9990 => x"72",
          9991 => x"74",
          9992 => x"4f",
          9993 => x"20",
          9994 => x"69",
          9995 => x"72",
          9996 => x"74",
          9997 => x"41",
          9998 => x"20",
          9999 => x"69",
         10000 => x"72",
         10001 => x"74",
         10002 => x"41",
         10003 => x"20",
         10004 => x"69",
         10005 => x"72",
         10006 => x"74",
         10007 => x"41",
         10008 => x"20",
         10009 => x"69",
         10010 => x"72",
         10011 => x"74",
         10012 => x"41",
         10013 => x"20",
         10014 => x"69",
         10015 => x"72",
         10016 => x"74",
         10017 => x"65",
         10018 => x"6e",
         10019 => x"70",
         10020 => x"6d",
         10021 => x"2e",
         10022 => x"6e",
         10023 => x"69",
         10024 => x"74",
         10025 => x"72",
         10026 => x"00",
         10027 => x"75",
         10028 => x"78",
         10029 => x"62",
         10030 => x"00",
         10031 => x"4f",
         10032 => x"73",
         10033 => x"3a",
         10034 => x"61",
         10035 => x"64",
         10036 => x"20",
         10037 => x"74",
         10038 => x"69",
         10039 => x"73",
         10040 => x"61",
         10041 => x"30",
         10042 => x"6c",
         10043 => x"65",
         10044 => x"69",
         10045 => x"61",
         10046 => x"6c",
         10047 => x"00",
         10048 => x"20",
         10049 => x"6c",
         10050 => x"69",
         10051 => x"2e",
         10052 => x"00",
         10053 => x"6f",
         10054 => x"6e",
         10055 => x"2e",
         10056 => x"6f",
         10057 => x"72",
         10058 => x"2e",
         10059 => x"00",
         10060 => x"30",
         10061 => x"28",
         10062 => x"78",
         10063 => x"25",
         10064 => x"78",
         10065 => x"38",
         10066 => x"00",
         10067 => x"75",
         10068 => x"4d",
         10069 => x"72",
         10070 => x"43",
         10071 => x"6c",
         10072 => x"2e",
         10073 => x"30",
         10074 => x"20",
         10075 => x"58",
         10076 => x"3f",
         10077 => x"30",
         10078 => x"20",
         10079 => x"58",
         10080 => x"30",
         10081 => x"20",
         10082 => x"6c",
         10083 => x"00",
         10084 => x"78",
         10085 => x"74",
         10086 => x"20",
         10087 => x"65",
         10088 => x"25",
         10089 => x"78",
         10090 => x"2e",
         10091 => x"61",
         10092 => x"6e",
         10093 => x"6f",
         10094 => x"40",
         10095 => x"38",
         10096 => x"2e",
         10097 => x"00",
         10098 => x"61",
         10099 => x"72",
         10100 => x"72",
         10101 => x"20",
         10102 => x"65",
         10103 => x"64",
         10104 => x"00",
         10105 => x"65",
         10106 => x"72",
         10107 => x"67",
         10108 => x"70",
         10109 => x"61",
         10110 => x"6e",
         10111 => x"00",
         10112 => x"6f",
         10113 => x"72",
         10114 => x"6f",
         10115 => x"67",
         10116 => x"00",
         10117 => x"50",
         10118 => x"69",
         10119 => x"64",
         10120 => x"73",
         10121 => x"2e",
         10122 => x"00",
         10123 => x"64",
         10124 => x"73",
         10125 => x"00",
         10126 => x"64",
         10127 => x"73",
         10128 => x"61",
         10129 => x"6f",
         10130 => x"6e",
         10131 => x"00",
         10132 => x"65",
         10133 => x"79",
         10134 => x"68",
         10135 => x"74",
         10136 => x"20",
         10137 => x"6e",
         10138 => x"70",
         10139 => x"65",
         10140 => x"63",
         10141 => x"61",
         10142 => x"00",
         10143 => x"65",
         10144 => x"6e",
         10145 => x"72",
         10146 => x"66",
         10147 => x"75",
         10148 => x"6e",
         10149 => x"2e",
         10150 => x"6e",
         10151 => x"69",
         10152 => x"69",
         10153 => x"72",
         10154 => x"74",
         10155 => x"2e",
         10156 => x"64",
         10157 => x"2f",
         10158 => x"25",
         10159 => x"64",
         10160 => x"2e",
         10161 => x"64",
         10162 => x"6f",
         10163 => x"6f",
         10164 => x"67",
         10165 => x"74",
         10166 => x"00",
         10167 => x"28",
         10168 => x"6d",
         10169 => x"43",
         10170 => x"6e",
         10171 => x"29",
         10172 => x"0a",
         10173 => x"69",
         10174 => x"20",
         10175 => x"6c",
         10176 => x"6e",
         10177 => x"3a",
         10178 => x"20",
         10179 => x"42",
         10180 => x"52",
         10181 => x"20",
         10182 => x"38",
         10183 => x"30",
         10184 => x"2e",
         10185 => x"20",
         10186 => x"44",
         10187 => x"20",
         10188 => x"20",
         10189 => x"38",
         10190 => x"30",
         10191 => x"2e",
         10192 => x"20",
         10193 => x"4e",
         10194 => x"42",
         10195 => x"20",
         10196 => x"38",
         10197 => x"30",
         10198 => x"2e",
         10199 => x"20",
         10200 => x"52",
         10201 => x"20",
         10202 => x"20",
         10203 => x"38",
         10204 => x"30",
         10205 => x"2e",
         10206 => x"20",
         10207 => x"41",
         10208 => x"20",
         10209 => x"20",
         10210 => x"38",
         10211 => x"30",
         10212 => x"2e",
         10213 => x"20",
         10214 => x"44",
         10215 => x"52",
         10216 => x"20",
         10217 => x"76",
         10218 => x"73",
         10219 => x"30",
         10220 => x"2e",
         10221 => x"20",
         10222 => x"49",
         10223 => x"31",
         10224 => x"20",
         10225 => x"6d",
         10226 => x"20",
         10227 => x"30",
         10228 => x"2e",
         10229 => x"20",
         10230 => x"4e",
         10231 => x"43",
         10232 => x"20",
         10233 => x"61",
         10234 => x"6c",
         10235 => x"30",
         10236 => x"2e",
         10237 => x"20",
         10238 => x"49",
         10239 => x"4f",
         10240 => x"42",
         10241 => x"00",
         10242 => x"20",
         10243 => x"42",
         10244 => x"43",
         10245 => x"20",
         10246 => x"4f",
         10247 => x"00",
         10248 => x"20",
         10249 => x"53",
         10250 => x"20",
         10251 => x"50",
         10252 => x"64",
         10253 => x"73",
         10254 => x"3a",
         10255 => x"20",
         10256 => x"50",
         10257 => x"65",
         10258 => x"20",
         10259 => x"74",
         10260 => x"41",
         10261 => x"65",
         10262 => x"3d",
         10263 => x"38",
         10264 => x"00",
         10265 => x"20",
         10266 => x"50",
         10267 => x"65",
         10268 => x"79",
         10269 => x"61",
         10270 => x"41",
         10271 => x"65",
         10272 => x"3d",
         10273 => x"38",
         10274 => x"00",
         10275 => x"20",
         10276 => x"74",
         10277 => x"20",
         10278 => x"72",
         10279 => x"64",
         10280 => x"73",
         10281 => x"20",
         10282 => x"3d",
         10283 => x"38",
         10284 => x"00",
         10285 => x"69",
         10286 => x"00",
         10287 => x"20",
         10288 => x"50",
         10289 => x"64",
         10290 => x"20",
         10291 => x"20",
         10292 => x"20",
         10293 => x"20",
         10294 => x"3d",
         10295 => x"34",
         10296 => x"00",
         10297 => x"20",
         10298 => x"79",
         10299 => x"6d",
         10300 => x"6f",
         10301 => x"46",
         10302 => x"20",
         10303 => x"20",
         10304 => x"3d",
         10305 => x"2e",
         10306 => x"64",
         10307 => x"0a",
         10308 => x"20",
         10309 => x"44",
         10310 => x"20",
         10311 => x"63",
         10312 => x"72",
         10313 => x"20",
         10314 => x"20",
         10315 => x"3d",
         10316 => x"2e",
         10317 => x"64",
         10318 => x"0a",
         10319 => x"20",
         10320 => x"69",
         10321 => x"6f",
         10322 => x"53",
         10323 => x"4d",
         10324 => x"6f",
         10325 => x"46",
         10326 => x"3d",
         10327 => x"2e",
         10328 => x"64",
         10329 => x"0a",
         10330 => x"6d",
         10331 => x"00",
         10332 => x"65",
         10333 => x"6d",
         10334 => x"6c",
         10335 => x"00",
         10336 => x"56",
         10337 => x"56",
         10338 => x"00",
         10339 => x"6e",
         10340 => x"77",
         10341 => x"00",
         10342 => x"00",
         10343 => x"00",
         10344 => x"00",
         10345 => x"00",
         10346 => x"00",
         10347 => x"00",
         10348 => x"00",
         10349 => x"00",
         10350 => x"00",
         10351 => x"00",
         10352 => x"00",
         10353 => x"00",
         10354 => x"00",
         10355 => x"00",
         10356 => x"00",
         10357 => x"00",
         10358 => x"00",
         10359 => x"00",
         10360 => x"00",
         10361 => x"00",
         10362 => x"00",
         10363 => x"00",
         10364 => x"00",
         10365 => x"00",
         10366 => x"00",
         10367 => x"00",
         10368 => x"00",
         10369 => x"00",
         10370 => x"00",
         10371 => x"00",
         10372 => x"00",
         10373 => x"00",
         10374 => x"00",
         10375 => x"00",
         10376 => x"00",
         10377 => x"00",
         10378 => x"00",
         10379 => x"00",
         10380 => x"00",
         10381 => x"00",
         10382 => x"00",
         10383 => x"00",
         10384 => x"00",
         10385 => x"00",
         10386 => x"00",
         10387 => x"00",
         10388 => x"00",
         10389 => x"00",
         10390 => x"00",
         10391 => x"00",
         10392 => x"00",
         10393 => x"00",
         10394 => x"00",
         10395 => x"00",
         10396 => x"00",
         10397 => x"00",
         10398 => x"00",
         10399 => x"00",
         10400 => x"00",
         10401 => x"00",
         10402 => x"00",
         10403 => x"00",
         10404 => x"00",
         10405 => x"00",
         10406 => x"00",
         10407 => x"5b",
         10408 => x"5b",
         10409 => x"5b",
         10410 => x"5b",
         10411 => x"5b",
         10412 => x"5b",
         10413 => x"5b",
         10414 => x"30",
         10415 => x"5b",
         10416 => x"5b",
         10417 => x"5b",
         10418 => x"00",
         10419 => x"00",
         10420 => x"00",
         10421 => x"00",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"69",
         10430 => x"72",
         10431 => x"69",
         10432 => x"00",
         10433 => x"00",
         10434 => x"30",
         10435 => x"20",
         10436 => x"0a",
         10437 => x"61",
         10438 => x"64",
         10439 => x"20",
         10440 => x"65",
         10441 => x"68",
         10442 => x"69",
         10443 => x"72",
         10444 => x"69",
         10445 => x"74",
         10446 => x"4f",
         10447 => x"00",
         10448 => x"61",
         10449 => x"74",
         10450 => x"65",
         10451 => x"72",
         10452 => x"65",
         10453 => x"73",
         10454 => x"79",
         10455 => x"6c",
         10456 => x"64",
         10457 => x"62",
         10458 => x"67",
         10459 => x"44",
         10460 => x"2a",
         10461 => x"3f",
         10462 => x"00",
         10463 => x"2c",
         10464 => x"5d",
         10465 => x"41",
         10466 => x"41",
         10467 => x"00",
         10468 => x"fe",
         10469 => x"44",
         10470 => x"2e",
         10471 => x"4f",
         10472 => x"4d",
         10473 => x"20",
         10474 => x"54",
         10475 => x"20",
         10476 => x"4f",
         10477 => x"4d",
         10478 => x"20",
         10479 => x"54",
         10480 => x"20",
         10481 => x"00",
         10482 => x"00",
         10483 => x"00",
         10484 => x"00",
         10485 => x"03",
         10486 => x"0e",
         10487 => x"16",
         10488 => x"00",
         10489 => x"9a",
         10490 => x"41",
         10491 => x"45",
         10492 => x"49",
         10493 => x"92",
         10494 => x"4f",
         10495 => x"99",
         10496 => x"9d",
         10497 => x"49",
         10498 => x"a5",
         10499 => x"a9",
         10500 => x"ad",
         10501 => x"b1",
         10502 => x"b5",
         10503 => x"b9",
         10504 => x"bd",
         10505 => x"c1",
         10506 => x"c5",
         10507 => x"c9",
         10508 => x"cd",
         10509 => x"d1",
         10510 => x"d5",
         10511 => x"d9",
         10512 => x"dd",
         10513 => x"e1",
         10514 => x"e5",
         10515 => x"e9",
         10516 => x"ed",
         10517 => x"f1",
         10518 => x"f5",
         10519 => x"f9",
         10520 => x"fd",
         10521 => x"2e",
         10522 => x"5b",
         10523 => x"22",
         10524 => x"3e",
         10525 => x"00",
         10526 => x"01",
         10527 => x"10",
         10528 => x"00",
         10529 => x"00",
         10530 => x"01",
         10531 => x"04",
         10532 => x"10",
         10533 => x"00",
         10534 => x"c7",
         10535 => x"e9",
         10536 => x"e4",
         10537 => x"e5",
         10538 => x"ea",
         10539 => x"e8",
         10540 => x"ee",
         10541 => x"c4",
         10542 => x"c9",
         10543 => x"c6",
         10544 => x"f6",
         10545 => x"fb",
         10546 => x"ff",
         10547 => x"dc",
         10548 => x"a3",
         10549 => x"a7",
         10550 => x"e1",
         10551 => x"f3",
         10552 => x"f1",
         10553 => x"aa",
         10554 => x"bf",
         10555 => x"ac",
         10556 => x"bc",
         10557 => x"ab",
         10558 => x"91",
         10559 => x"93",
         10560 => x"24",
         10561 => x"62",
         10562 => x"55",
         10563 => x"51",
         10564 => x"5d",
         10565 => x"5b",
         10566 => x"14",
         10567 => x"2c",
         10568 => x"00",
         10569 => x"5e",
         10570 => x"5a",
         10571 => x"69",
         10572 => x"60",
         10573 => x"6c",
         10574 => x"68",
         10575 => x"65",
         10576 => x"58",
         10577 => x"53",
         10578 => x"6a",
         10579 => x"0c",
         10580 => x"84",
         10581 => x"90",
         10582 => x"b1",
         10583 => x"93",
         10584 => x"a3",
         10585 => x"b5",
         10586 => x"a6",
         10587 => x"a9",
         10588 => x"1e",
         10589 => x"b5",
         10590 => x"61",
         10591 => x"65",
         10592 => x"20",
         10593 => x"f7",
         10594 => x"b0",
         10595 => x"b7",
         10596 => x"7f",
         10597 => x"a0",
         10598 => x"61",
         10599 => x"e0",
         10600 => x"f8",
         10601 => x"ff",
         10602 => x"78",
         10603 => x"30",
         10604 => x"06",
         10605 => x"10",
         10606 => x"2e",
         10607 => x"06",
         10608 => x"4d",
         10609 => x"81",
         10610 => x"82",
         10611 => x"84",
         10612 => x"87",
         10613 => x"89",
         10614 => x"8b",
         10615 => x"8d",
         10616 => x"8f",
         10617 => x"91",
         10618 => x"93",
         10619 => x"f6",
         10620 => x"97",
         10621 => x"98",
         10622 => x"9b",
         10623 => x"9d",
         10624 => x"9f",
         10625 => x"a0",
         10626 => x"a2",
         10627 => x"a4",
         10628 => x"a7",
         10629 => x"a9",
         10630 => x"ab",
         10631 => x"ac",
         10632 => x"af",
         10633 => x"b1",
         10634 => x"b3",
         10635 => x"b5",
         10636 => x"b7",
         10637 => x"b8",
         10638 => x"bb",
         10639 => x"bc",
         10640 => x"f7",
         10641 => x"c1",
         10642 => x"c3",
         10643 => x"c5",
         10644 => x"c7",
         10645 => x"c7",
         10646 => x"cb",
         10647 => x"cd",
         10648 => x"dd",
         10649 => x"8e",
         10650 => x"12",
         10651 => x"03",
         10652 => x"f4",
         10653 => x"f8",
         10654 => x"22",
         10655 => x"3a",
         10656 => x"65",
         10657 => x"3b",
         10658 => x"66",
         10659 => x"40",
         10660 => x"41",
         10661 => x"0a",
         10662 => x"40",
         10663 => x"86",
         10664 => x"89",
         10665 => x"58",
         10666 => x"5a",
         10667 => x"5c",
         10668 => x"5e",
         10669 => x"93",
         10670 => x"62",
         10671 => x"64",
         10672 => x"66",
         10673 => x"97",
         10674 => x"6a",
         10675 => x"6c",
         10676 => x"6e",
         10677 => x"70",
         10678 => x"9d",
         10679 => x"74",
         10680 => x"76",
         10681 => x"78",
         10682 => x"7a",
         10683 => x"7c",
         10684 => x"7e",
         10685 => x"a6",
         10686 => x"82",
         10687 => x"84",
         10688 => x"86",
         10689 => x"ae",
         10690 => x"b1",
         10691 => x"45",
         10692 => x"8e",
         10693 => x"90",
         10694 => x"b7",
         10695 => x"03",
         10696 => x"fe",
         10697 => x"ac",
         10698 => x"86",
         10699 => x"89",
         10700 => x"b1",
         10701 => x"c2",
         10702 => x"a3",
         10703 => x"c4",
         10704 => x"cc",
         10705 => x"8c",
         10706 => x"8f",
         10707 => x"18",
         10708 => x"0a",
         10709 => x"f3",
         10710 => x"f5",
         10711 => x"f7",
         10712 => x"f9",
         10713 => x"fa",
         10714 => x"20",
         10715 => x"10",
         10716 => x"22",
         10717 => x"36",
         10718 => x"0e",
         10719 => x"01",
         10720 => x"d0",
         10721 => x"61",
         10722 => x"00",
         10723 => x"7d",
         10724 => x"63",
         10725 => x"96",
         10726 => x"5a",
         10727 => x"08",
         10728 => x"06",
         10729 => x"08",
         10730 => x"08",
         10731 => x"06",
         10732 => x"07",
         10733 => x"52",
         10734 => x"54",
         10735 => x"56",
         10736 => x"60",
         10737 => x"70",
         10738 => x"ba",
         10739 => x"c8",
         10740 => x"ca",
         10741 => x"da",
         10742 => x"f8",
         10743 => x"ea",
         10744 => x"fa",
         10745 => x"80",
         10746 => x"90",
         10747 => x"a0",
         10748 => x"b0",
         10749 => x"b8",
         10750 => x"b2",
         10751 => x"cc",
         10752 => x"c3",
         10753 => x"02",
         10754 => x"02",
         10755 => x"01",
         10756 => x"f3",
         10757 => x"fc",
         10758 => x"01",
         10759 => x"70",
         10760 => x"84",
         10761 => x"83",
         10762 => x"1a",
         10763 => x"2f",
         10764 => x"02",
         10765 => x"06",
         10766 => x"02",
         10767 => x"64",
         10768 => x"26",
         10769 => x"1a",
         10770 => x"00",
         10771 => x"00",
         10772 => x"02",
         10773 => x"00",
         10774 => x"00",
         10775 => x"00",
         10776 => x"04",
         10777 => x"00",
         10778 => x"00",
         10779 => x"00",
         10780 => x"14",
         10781 => x"00",
         10782 => x"00",
         10783 => x"00",
         10784 => x"2b",
         10785 => x"00",
         10786 => x"00",
         10787 => x"00",
         10788 => x"30",
         10789 => x"00",
         10790 => x"00",
         10791 => x"00",
         10792 => x"3c",
         10793 => x"00",
         10794 => x"00",
         10795 => x"00",
         10796 => x"3d",
         10797 => x"00",
         10798 => x"00",
         10799 => x"00",
         10800 => x"3f",
         10801 => x"00",
         10802 => x"00",
         10803 => x"00",
         10804 => x"40",
         10805 => x"00",
         10806 => x"00",
         10807 => x"00",
         10808 => x"41",
         10809 => x"00",
         10810 => x"00",
         10811 => x"00",
         10812 => x"42",
         10813 => x"00",
         10814 => x"00",
         10815 => x"00",
         10816 => x"43",
         10817 => x"00",
         10818 => x"00",
         10819 => x"00",
         10820 => x"50",
         10821 => x"00",
         10822 => x"00",
         10823 => x"00",
         10824 => x"51",
         10825 => x"00",
         10826 => x"00",
         10827 => x"00",
         10828 => x"54",
         10829 => x"00",
         10830 => x"00",
         10831 => x"00",
         10832 => x"55",
         10833 => x"00",
         10834 => x"00",
         10835 => x"00",
         10836 => x"79",
         10837 => x"00",
         10838 => x"00",
         10839 => x"00",
         10840 => x"78",
         10841 => x"00",
         10842 => x"00",
         10843 => x"00",
         10844 => x"82",
         10845 => x"00",
         10846 => x"00",
         10847 => x"00",
         10848 => x"83",
         10849 => x"00",
         10850 => x"00",
         10851 => x"00",
         10852 => x"85",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"87",
         10857 => x"00",
         10858 => x"00",
         10859 => x"00",
         10860 => x"8c",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"8d",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"8e",
         10869 => x"00",
         10870 => x"00",
         10871 => x"00",
         10872 => x"8f",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"01",
         10881 => x"00",
         10882 => x"01",
         10883 => x"81",
         10884 => x"00",
         10885 => x"7f",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"f5",
         10891 => x"f5",
         10892 => x"f5",
         10893 => x"00",
         10894 => x"01",
         10895 => x"01",
         10896 => x"01",
         10897 => x"00",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"00",
         10927 => x"00",
         10928 => x"e0",
         10929 => x"cf",
         10930 => x"f9",
         10931 => x"fd",
         10932 => x"c1",
         10933 => x"c5",
         10934 => x"e4",
         10935 => x"ee",
         10936 => x"61",
         10937 => x"65",
         10938 => x"69",
         10939 => x"2a",
         10940 => x"21",
         10941 => x"25",
         10942 => x"29",
         10943 => x"2b",
         10944 => x"01",
         10945 => x"05",
         10946 => x"09",
         10947 => x"0d",
         10948 => x"11",
         10949 => x"15",
         10950 => x"19",
         10951 => x"54",
         10952 => x"81",
         10953 => x"85",
         10954 => x"89",
         10955 => x"8d",
         10956 => x"91",
         10957 => x"95",
         10958 => x"99",
         10959 => x"40",
         10960 => x"e8",
         10961 => x"00",
         10962 => x"00",
         10963 => x"00",
         10964 => x"00",
         10965 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"cc",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"9f",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"8b",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"84",
           393 => x"82",
           394 => x"af",
           395 => x"d6",
           396 => x"80",
           397 => x"d6",
           398 => x"ad",
           399 => x"e4",
           400 => x"90",
           401 => x"e4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"84",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"84",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"84",
           416 => x"82",
           417 => x"93",
           418 => x"d6",
           419 => x"80",
           420 => x"d6",
           421 => x"c0",
           422 => x"e4",
           423 => x"90",
           424 => x"e4",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"f0",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"d6",
           636 => x"05",
           637 => x"e4",
           638 => x"08",
           639 => x"e4",
           640 => x"08",
           641 => x"bc",
           642 => x"84",
           643 => x"d6",
           644 => x"82",
           645 => x"f8",
           646 => x"d6",
           647 => x"05",
           648 => x"d6",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"e4",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"e4",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"e4",
           668 => x"08",
           669 => x"d6",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"d6",
           674 => x"05",
           675 => x"e4",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"d6",
           681 => x"05",
           682 => x"e9",
           683 => x"e4",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"e4",
           688 => x"0c",
           689 => x"e4",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"e4",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"d6",
           698 => x"05",
           699 => x"71",
           700 => x"d6",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"d6",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"e4",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"d6",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"e4",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"e4",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"d6",
           736 => x"05",
           737 => x"d6",
           738 => x"05",
           739 => x"d6",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"d6",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"e4",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"d6",
           763 => x"05",
           764 => x"d6",
           765 => x"05",
           766 => x"d6",
           767 => x"05",
           768 => x"a3",
           769 => x"d8",
           770 => x"d6",
           771 => x"05",
           772 => x"e4",
           773 => x"08",
           774 => x"d8",
           775 => x"87",
           776 => x"d6",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"e4",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"e4",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"d6",
           797 => x"05",
           798 => x"33",
           799 => x"d6",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"e4",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"d6",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"d6",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"d6",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"e4",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"d6",
           856 => x"05",
           857 => x"e4",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"e4",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"e4",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"e4",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"e4",
           894 => x"0c",
           895 => x"e4",
           896 => x"08",
           897 => x"92",
           898 => x"d6",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"e4",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"e4",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"e4",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"e4",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"e4",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"e4",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"d6",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"d6",
           960 => x"05",
           961 => x"51",
           962 => x"d6",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"e4",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"d6",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"e4",
           983 => x"08",
           984 => x"83",
           985 => x"d8",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"e4",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"e4",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"d6",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"e4",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"d6",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"d6",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"d6",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"d6",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"d6",
          1055 => x"05",
          1056 => x"e4",
          1057 => x"08",
          1058 => x"d6",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"d6",
          1065 => x"05",
          1066 => x"e4",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"e4",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"e4",
          1082 => x"23",
          1083 => x"88",
          1084 => x"e4",
          1085 => x"23",
          1086 => x"d6",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"d6",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"d6",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"d6",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"d6",
          1111 => x"05",
          1112 => x"e4",
          1113 => x"08",
          1114 => x"d6",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"d6",
          1121 => x"05",
          1122 => x"e4",
          1123 => x"22",
          1124 => x"51",
          1125 => x"d6",
          1126 => x"05",
          1127 => x"e8",
          1128 => x"e4",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"d6",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"d6",
          1142 => x"05",
          1143 => x"e4",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"e4",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"d6",
          1162 => x"05",
          1163 => x"d6",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"e4",
          1177 => x"0c",
          1178 => x"e4",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"d6",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"e4",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"d6",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"d6",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"d6",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"d6",
          1224 => x"05",
          1225 => x"e4",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"e4",
          1235 => x"33",
          1236 => x"70",
          1237 => x"d6",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"d6",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"e4",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"e4",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"e4",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"d6",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"e4",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"d6",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"d6",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"d6",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"d6",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"e4",
          1382 => x"22",
          1383 => x"54",
          1384 => x"e4",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"e4",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"e4",
          1398 => x"08",
          1399 => x"e4",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"e4",
          1408 => x"22",
          1409 => x"53",
          1410 => x"e4",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"d6",
          1416 => x"05",
          1417 => x"d6",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"e4",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"e4",
          1431 => x"22",
          1432 => x"53",
          1433 => x"e4",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"d6",
          1439 => x"05",
          1440 => x"d6",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"e4",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"d6",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"e4",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"d6",
          1468 => x"05",
          1469 => x"54",
          1470 => x"d6",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"d6",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"e4",
          1480 => x"08",
          1481 => x"e4",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"d6",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"d6",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"e4",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"e4",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"e4",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"e4",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"e4",
          1521 => x"08",
          1522 => x"e4",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"d8",
          1527 => x"3d",
          1528 => x"e4",
          1529 => x"d6",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"e4",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"e4",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"f2",
          1556 => x"f2",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"d6",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"bc",
          1568 => x"bc",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"d6",
          1577 => x"05",
          1578 => x"d6",
          1579 => x"05",
          1580 => x"d6",
          1581 => x"05",
          1582 => x"d8",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"e4",
          1586 => x"d6",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"d6",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"e4",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"e4",
          1604 => x"08",
          1605 => x"d6",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"d6",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"e4",
          1626 => x"08",
          1627 => x"e4",
          1628 => x"0c",
          1629 => x"e4",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"e4",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"e4",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"e4",
          1646 => x"d6",
          1647 => x"3d",
          1648 => x"e4",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"d6",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"e4",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"d6",
          1683 => x"05",
          1684 => x"d6",
          1685 => x"05",
          1686 => x"80",
          1687 => x"d6",
          1688 => x"05",
          1689 => x"e4",
          1690 => x"08",
          1691 => x"e4",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"d8",
          1697 => x"a3",
          1698 => x"e4",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"e4",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"d6",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"d6",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"d6",
          1733 => x"05",
          1734 => x"e4",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"d6",
          1744 => x"05",
          1745 => x"33",
          1746 => x"e4",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"d6",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"e4",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"e4",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"d6",
          1778 => x"05",
          1779 => x"e4",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"e4",
          1785 => x"0c",
          1786 => x"e4",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"e4",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"e4",
          1796 => x"0c",
          1797 => x"e4",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"d6",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"d6",
          1809 => x"05",
          1810 => x"e4",
          1811 => x"08",
          1812 => x"e4",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"e4",
          1816 => x"0c",
          1817 => x"d6",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"e4",
          1822 => x"08",
          1823 => x"06",
          1824 => x"e4",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"d6",
          1829 => x"3d",
          1830 => x"e4",
          1831 => x"d6",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"d6",
          1835 => x"05",
          1836 => x"e4",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"d6",
          1842 => x"05",
          1843 => x"82",
          1844 => x"d6",
          1845 => x"05",
          1846 => x"e4",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"d6",
          1862 => x"05",
          1863 => x"e4",
          1864 => x"08",
          1865 => x"e4",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"e4",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"e4",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"e4",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"e4",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"d6",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"e4",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"e4",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"e4",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"d6",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"e4",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"e4",
          1939 => x"08",
          1940 => x"d6",
          1941 => x"05",
          1942 => x"e4",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"d8",
          1947 => x"3d",
          1948 => x"e4",
          1949 => x"d6",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"d6",
          1953 => x"05",
          1954 => x"e4",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"d6",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"d6",
          1963 => x"05",
          1964 => x"70",
          1965 => x"d6",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"e4",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"d6",
          1985 => x"05",
          1986 => x"e4",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"e4",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"e4",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"e4",
          2005 => x"08",
          2006 => x"d6",
          2007 => x"05",
          2008 => x"e4",
          2009 => x"08",
          2010 => x"71",
          2011 => x"e4",
          2012 => x"08",
          2013 => x"d6",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"e4",
          2022 => x"d6",
          2023 => x"3d",
          2024 => x"e4",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"e4",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"d6",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"e4",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"e4",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"e4",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"e4",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"e4",
          2082 => x"08",
          2083 => x"71",
          2084 => x"d6",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"d6",
          2089 => x"05",
          2090 => x"e4",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"e4",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"52",
          2100 => x"08",
          2101 => x"51",
          2102 => x"82",
          2103 => x"70",
          2104 => x"08",
          2105 => x"82",
          2106 => x"f8",
          2107 => x"05",
          2108 => x"54",
          2109 => x"3f",
          2110 => x"08",
          2111 => x"e4",
          2112 => x"0c",
          2113 => x"e4",
          2114 => x"08",
          2115 => x"0b",
          2116 => x"08",
          2117 => x"bc",
          2118 => x"e4",
          2119 => x"08",
          2120 => x"08",
          2121 => x"05",
          2122 => x"34",
          2123 => x"08",
          2124 => x"53",
          2125 => x"08",
          2126 => x"52",
          2127 => x"08",
          2128 => x"51",
          2129 => x"82",
          2130 => x"70",
          2131 => x"08",
          2132 => x"54",
          2133 => x"08",
          2134 => x"82",
          2135 => x"88",
          2136 => x"d6",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"d6",
          2143 => x"05",
          2144 => x"e4",
          2145 => x"08",
          2146 => x"0b",
          2147 => x"08",
          2148 => x"80",
          2149 => x"d6",
          2150 => x"05",
          2151 => x"33",
          2152 => x"08",
          2153 => x"81",
          2154 => x"e4",
          2155 => x"0c",
          2156 => x"06",
          2157 => x"80",
          2158 => x"82",
          2159 => x"8c",
          2160 => x"05",
          2161 => x"08",
          2162 => x"82",
          2163 => x"8c",
          2164 => x"2e",
          2165 => x"be",
          2166 => x"e4",
          2167 => x"08",
          2168 => x"d6",
          2169 => x"05",
          2170 => x"e4",
          2171 => x"08",
          2172 => x"08",
          2173 => x"31",
          2174 => x"e4",
          2175 => x"0c",
          2176 => x"e4",
          2177 => x"08",
          2178 => x"0c",
          2179 => x"82",
          2180 => x"04",
          2181 => x"08",
          2182 => x"e4",
          2183 => x"0d",
          2184 => x"08",
          2185 => x"82",
          2186 => x"fc",
          2187 => x"d6",
          2188 => x"05",
          2189 => x"80",
          2190 => x"d6",
          2191 => x"05",
          2192 => x"82",
          2193 => x"90",
          2194 => x"d6",
          2195 => x"05",
          2196 => x"82",
          2197 => x"90",
          2198 => x"d6",
          2199 => x"05",
          2200 => x"a9",
          2201 => x"e4",
          2202 => x"08",
          2203 => x"d6",
          2204 => x"05",
          2205 => x"71",
          2206 => x"d6",
          2207 => x"05",
          2208 => x"82",
          2209 => x"fc",
          2210 => x"be",
          2211 => x"e4",
          2212 => x"08",
          2213 => x"d8",
          2214 => x"3d",
          2215 => x"e4",
          2216 => x"d6",
          2217 => x"82",
          2218 => x"f9",
          2219 => x"0b",
          2220 => x"08",
          2221 => x"82",
          2222 => x"88",
          2223 => x"25",
          2224 => x"d6",
          2225 => x"05",
          2226 => x"d6",
          2227 => x"05",
          2228 => x"82",
          2229 => x"f4",
          2230 => x"d6",
          2231 => x"05",
          2232 => x"81",
          2233 => x"e4",
          2234 => x"0c",
          2235 => x"08",
          2236 => x"82",
          2237 => x"fc",
          2238 => x"d6",
          2239 => x"05",
          2240 => x"b9",
          2241 => x"e4",
          2242 => x"08",
          2243 => x"e4",
          2244 => x"0c",
          2245 => x"d6",
          2246 => x"05",
          2247 => x"e4",
          2248 => x"08",
          2249 => x"0b",
          2250 => x"08",
          2251 => x"82",
          2252 => x"f0",
          2253 => x"d6",
          2254 => x"05",
          2255 => x"82",
          2256 => x"8c",
          2257 => x"82",
          2258 => x"88",
          2259 => x"82",
          2260 => x"d6",
          2261 => x"82",
          2262 => x"f8",
          2263 => x"82",
          2264 => x"fc",
          2265 => x"2e",
          2266 => x"d6",
          2267 => x"05",
          2268 => x"d6",
          2269 => x"05",
          2270 => x"e4",
          2271 => x"08",
          2272 => x"d8",
          2273 => x"3d",
          2274 => x"e4",
          2275 => x"d6",
          2276 => x"82",
          2277 => x"fb",
          2278 => x"0b",
          2279 => x"08",
          2280 => x"82",
          2281 => x"88",
          2282 => x"25",
          2283 => x"d6",
          2284 => x"05",
          2285 => x"d6",
          2286 => x"05",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"d6",
          2290 => x"05",
          2291 => x"90",
          2292 => x"e4",
          2293 => x"08",
          2294 => x"e4",
          2295 => x"0c",
          2296 => x"d6",
          2297 => x"05",
          2298 => x"d6",
          2299 => x"05",
          2300 => x"a2",
          2301 => x"d8",
          2302 => x"d6",
          2303 => x"05",
          2304 => x"d6",
          2305 => x"05",
          2306 => x"90",
          2307 => x"e4",
          2308 => x"08",
          2309 => x"e4",
          2310 => x"0c",
          2311 => x"08",
          2312 => x"70",
          2313 => x"0c",
          2314 => x"0d",
          2315 => x"0c",
          2316 => x"e4",
          2317 => x"d6",
          2318 => x"3d",
          2319 => x"82",
          2320 => x"8c",
          2321 => x"82",
          2322 => x"88",
          2323 => x"80",
          2324 => x"d6",
          2325 => x"82",
          2326 => x"54",
          2327 => x"82",
          2328 => x"04",
          2329 => x"08",
          2330 => x"e4",
          2331 => x"0d",
          2332 => x"d6",
          2333 => x"05",
          2334 => x"d6",
          2335 => x"05",
          2336 => x"3f",
          2337 => x"08",
          2338 => x"d8",
          2339 => x"3d",
          2340 => x"e4",
          2341 => x"d6",
          2342 => x"82",
          2343 => x"fd",
          2344 => x"0b",
          2345 => x"08",
          2346 => x"80",
          2347 => x"e4",
          2348 => x"0c",
          2349 => x"08",
          2350 => x"82",
          2351 => x"88",
          2352 => x"b9",
          2353 => x"e4",
          2354 => x"08",
          2355 => x"38",
          2356 => x"d6",
          2357 => x"05",
          2358 => x"38",
          2359 => x"08",
          2360 => x"10",
          2361 => x"08",
          2362 => x"82",
          2363 => x"fc",
          2364 => x"82",
          2365 => x"fc",
          2366 => x"b8",
          2367 => x"e4",
          2368 => x"08",
          2369 => x"e1",
          2370 => x"e4",
          2371 => x"08",
          2372 => x"08",
          2373 => x"26",
          2374 => x"d6",
          2375 => x"05",
          2376 => x"e4",
          2377 => x"08",
          2378 => x"e4",
          2379 => x"0c",
          2380 => x"08",
          2381 => x"82",
          2382 => x"fc",
          2383 => x"82",
          2384 => x"f8",
          2385 => x"d6",
          2386 => x"05",
          2387 => x"82",
          2388 => x"fc",
          2389 => x"d6",
          2390 => x"05",
          2391 => x"82",
          2392 => x"8c",
          2393 => x"95",
          2394 => x"e4",
          2395 => x"08",
          2396 => x"38",
          2397 => x"08",
          2398 => x"70",
          2399 => x"08",
          2400 => x"51",
          2401 => x"d6",
          2402 => x"05",
          2403 => x"d6",
          2404 => x"05",
          2405 => x"d6",
          2406 => x"05",
          2407 => x"d8",
          2408 => x"0d",
          2409 => x"0c",
          2410 => x"e4",
          2411 => x"d6",
          2412 => x"3d",
          2413 => x"82",
          2414 => x"f0",
          2415 => x"d6",
          2416 => x"05",
          2417 => x"73",
          2418 => x"e4",
          2419 => x"08",
          2420 => x"53",
          2421 => x"72",
          2422 => x"08",
          2423 => x"72",
          2424 => x"53",
          2425 => x"09",
          2426 => x"38",
          2427 => x"08",
          2428 => x"70",
          2429 => x"71",
          2430 => x"39",
          2431 => x"08",
          2432 => x"53",
          2433 => x"09",
          2434 => x"38",
          2435 => x"d6",
          2436 => x"05",
          2437 => x"e4",
          2438 => x"08",
          2439 => x"05",
          2440 => x"08",
          2441 => x"33",
          2442 => x"08",
          2443 => x"82",
          2444 => x"f8",
          2445 => x"72",
          2446 => x"81",
          2447 => x"38",
          2448 => x"08",
          2449 => x"70",
          2450 => x"71",
          2451 => x"51",
          2452 => x"82",
          2453 => x"f8",
          2454 => x"d6",
          2455 => x"05",
          2456 => x"e4",
          2457 => x"0c",
          2458 => x"08",
          2459 => x"80",
          2460 => x"38",
          2461 => x"08",
          2462 => x"80",
          2463 => x"38",
          2464 => x"90",
          2465 => x"e4",
          2466 => x"34",
          2467 => x"08",
          2468 => x"70",
          2469 => x"71",
          2470 => x"51",
          2471 => x"82",
          2472 => x"f8",
          2473 => x"a4",
          2474 => x"82",
          2475 => x"f4",
          2476 => x"d6",
          2477 => x"05",
          2478 => x"81",
          2479 => x"70",
          2480 => x"72",
          2481 => x"e4",
          2482 => x"34",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"72",
          2486 => x"38",
          2487 => x"d6",
          2488 => x"05",
          2489 => x"39",
          2490 => x"08",
          2491 => x"53",
          2492 => x"90",
          2493 => x"e4",
          2494 => x"33",
          2495 => x"26",
          2496 => x"39",
          2497 => x"d6",
          2498 => x"05",
          2499 => x"39",
          2500 => x"d6",
          2501 => x"05",
          2502 => x"82",
          2503 => x"f8",
          2504 => x"af",
          2505 => x"38",
          2506 => x"08",
          2507 => x"53",
          2508 => x"83",
          2509 => x"80",
          2510 => x"e4",
          2511 => x"0c",
          2512 => x"8a",
          2513 => x"e4",
          2514 => x"34",
          2515 => x"d6",
          2516 => x"05",
          2517 => x"e4",
          2518 => x"33",
          2519 => x"27",
          2520 => x"82",
          2521 => x"f8",
          2522 => x"80",
          2523 => x"94",
          2524 => x"e4",
          2525 => x"33",
          2526 => x"53",
          2527 => x"e4",
          2528 => x"34",
          2529 => x"08",
          2530 => x"d0",
          2531 => x"72",
          2532 => x"08",
          2533 => x"82",
          2534 => x"f8",
          2535 => x"90",
          2536 => x"38",
          2537 => x"08",
          2538 => x"f9",
          2539 => x"72",
          2540 => x"08",
          2541 => x"82",
          2542 => x"f8",
          2543 => x"72",
          2544 => x"38",
          2545 => x"d6",
          2546 => x"05",
          2547 => x"39",
          2548 => x"08",
          2549 => x"82",
          2550 => x"f4",
          2551 => x"54",
          2552 => x"8d",
          2553 => x"82",
          2554 => x"ec",
          2555 => x"f7",
          2556 => x"e4",
          2557 => x"33",
          2558 => x"e4",
          2559 => x"08",
          2560 => x"e4",
          2561 => x"33",
          2562 => x"d6",
          2563 => x"05",
          2564 => x"e4",
          2565 => x"08",
          2566 => x"05",
          2567 => x"08",
          2568 => x"55",
          2569 => x"82",
          2570 => x"f8",
          2571 => x"a5",
          2572 => x"e4",
          2573 => x"33",
          2574 => x"2e",
          2575 => x"d6",
          2576 => x"05",
          2577 => x"d6",
          2578 => x"05",
          2579 => x"e4",
          2580 => x"08",
          2581 => x"08",
          2582 => x"71",
          2583 => x"0b",
          2584 => x"08",
          2585 => x"82",
          2586 => x"ec",
          2587 => x"d6",
          2588 => x"3d",
          2589 => x"e4",
          2590 => x"d6",
          2591 => x"82",
          2592 => x"f7",
          2593 => x"0b",
          2594 => x"08",
          2595 => x"82",
          2596 => x"8c",
          2597 => x"80",
          2598 => x"d6",
          2599 => x"05",
          2600 => x"51",
          2601 => x"53",
          2602 => x"e4",
          2603 => x"34",
          2604 => x"06",
          2605 => x"2e",
          2606 => x"91",
          2607 => x"e4",
          2608 => x"08",
          2609 => x"05",
          2610 => x"ce",
          2611 => x"e4",
          2612 => x"33",
          2613 => x"2e",
          2614 => x"a4",
          2615 => x"82",
          2616 => x"f0",
          2617 => x"d6",
          2618 => x"05",
          2619 => x"81",
          2620 => x"70",
          2621 => x"72",
          2622 => x"e4",
          2623 => x"34",
          2624 => x"08",
          2625 => x"53",
          2626 => x"09",
          2627 => x"dc",
          2628 => x"e4",
          2629 => x"08",
          2630 => x"05",
          2631 => x"08",
          2632 => x"33",
          2633 => x"08",
          2634 => x"82",
          2635 => x"f8",
          2636 => x"d6",
          2637 => x"05",
          2638 => x"e4",
          2639 => x"08",
          2640 => x"b6",
          2641 => x"e4",
          2642 => x"08",
          2643 => x"84",
          2644 => x"39",
          2645 => x"d6",
          2646 => x"05",
          2647 => x"e4",
          2648 => x"08",
          2649 => x"05",
          2650 => x"08",
          2651 => x"33",
          2652 => x"08",
          2653 => x"81",
          2654 => x"0b",
          2655 => x"08",
          2656 => x"82",
          2657 => x"88",
          2658 => x"08",
          2659 => x"0c",
          2660 => x"53",
          2661 => x"d6",
          2662 => x"05",
          2663 => x"39",
          2664 => x"08",
          2665 => x"53",
          2666 => x"8d",
          2667 => x"82",
          2668 => x"ec",
          2669 => x"80",
          2670 => x"e4",
          2671 => x"33",
          2672 => x"27",
          2673 => x"d6",
          2674 => x"05",
          2675 => x"b9",
          2676 => x"8d",
          2677 => x"82",
          2678 => x"ec",
          2679 => x"d8",
          2680 => x"82",
          2681 => x"f4",
          2682 => x"39",
          2683 => x"08",
          2684 => x"53",
          2685 => x"90",
          2686 => x"e4",
          2687 => x"33",
          2688 => x"26",
          2689 => x"39",
          2690 => x"d6",
          2691 => x"05",
          2692 => x"39",
          2693 => x"d6",
          2694 => x"05",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"d6",
          2698 => x"05",
          2699 => x"73",
          2700 => x"38",
          2701 => x"08",
          2702 => x"53",
          2703 => x"27",
          2704 => x"d6",
          2705 => x"05",
          2706 => x"51",
          2707 => x"d6",
          2708 => x"05",
          2709 => x"e4",
          2710 => x"33",
          2711 => x"53",
          2712 => x"e4",
          2713 => x"34",
          2714 => x"08",
          2715 => x"53",
          2716 => x"ad",
          2717 => x"e4",
          2718 => x"33",
          2719 => x"53",
          2720 => x"e4",
          2721 => x"34",
          2722 => x"08",
          2723 => x"53",
          2724 => x"8d",
          2725 => x"82",
          2726 => x"ec",
          2727 => x"98",
          2728 => x"e4",
          2729 => x"33",
          2730 => x"08",
          2731 => x"54",
          2732 => x"26",
          2733 => x"0b",
          2734 => x"08",
          2735 => x"80",
          2736 => x"d6",
          2737 => x"05",
          2738 => x"d6",
          2739 => x"05",
          2740 => x"d6",
          2741 => x"05",
          2742 => x"82",
          2743 => x"fc",
          2744 => x"d6",
          2745 => x"05",
          2746 => x"81",
          2747 => x"70",
          2748 => x"52",
          2749 => x"33",
          2750 => x"08",
          2751 => x"fe",
          2752 => x"d6",
          2753 => x"05",
          2754 => x"80",
          2755 => x"82",
          2756 => x"fc",
          2757 => x"82",
          2758 => x"fc",
          2759 => x"d6",
          2760 => x"05",
          2761 => x"e4",
          2762 => x"08",
          2763 => x"81",
          2764 => x"e4",
          2765 => x"0c",
          2766 => x"08",
          2767 => x"82",
          2768 => x"8b",
          2769 => x"d6",
          2770 => x"f8",
          2771 => x"70",
          2772 => x"56",
          2773 => x"2e",
          2774 => x"8c",
          2775 => x"79",
          2776 => x"33",
          2777 => x"39",
          2778 => x"73",
          2779 => x"81",
          2780 => x"81",
          2781 => x"39",
          2782 => x"90",
          2783 => x"cc",
          2784 => x"52",
          2785 => x"3f",
          2786 => x"08",
          2787 => x"08",
          2788 => x"76",
          2789 => x"e7",
          2790 => x"d6",
          2791 => x"38",
          2792 => x"54",
          2793 => x"ff",
          2794 => x"17",
          2795 => x"06",
          2796 => x"77",
          2797 => x"ff",
          2798 => x"d6",
          2799 => x"3d",
          2800 => x"3d",
          2801 => x"71",
          2802 => x"8e",
          2803 => x"29",
          2804 => x"05",
          2805 => x"04",
          2806 => x"51",
          2807 => x"82",
          2808 => x"80",
          2809 => x"b2",
          2810 => x"f2",
          2811 => x"f8",
          2812 => x"39",
          2813 => x"51",
          2814 => x"82",
          2815 => x"80",
          2816 => x"b3",
          2817 => x"d6",
          2818 => x"bc",
          2819 => x"39",
          2820 => x"51",
          2821 => x"82",
          2822 => x"80",
          2823 => x"b4",
          2824 => x"39",
          2825 => x"51",
          2826 => x"b4",
          2827 => x"39",
          2828 => x"51",
          2829 => x"b4",
          2830 => x"39",
          2831 => x"51",
          2832 => x"b5",
          2833 => x"39",
          2834 => x"51",
          2835 => x"b5",
          2836 => x"39",
          2837 => x"51",
          2838 => x"b5",
          2839 => x"86",
          2840 => x"0d",
          2841 => x"0d",
          2842 => x"56",
          2843 => x"26",
          2844 => x"52",
          2845 => x"29",
          2846 => x"87",
          2847 => x"51",
          2848 => x"82",
          2849 => x"52",
          2850 => x"a5",
          2851 => x"d8",
          2852 => x"53",
          2853 => x"b6",
          2854 => x"ba",
          2855 => x"3d",
          2856 => x"3d",
          2857 => x"84",
          2858 => x"05",
          2859 => x"80",
          2860 => x"70",
          2861 => x"25",
          2862 => x"59",
          2863 => x"87",
          2864 => x"38",
          2865 => x"76",
          2866 => x"ff",
          2867 => x"93",
          2868 => x"82",
          2869 => x"76",
          2870 => x"70",
          2871 => x"92",
          2872 => x"d6",
          2873 => x"82",
          2874 => x"b9",
          2875 => x"d8",
          2876 => x"98",
          2877 => x"d6",
          2878 => x"96",
          2879 => x"54",
          2880 => x"77",
          2881 => x"81",
          2882 => x"82",
          2883 => x"57",
          2884 => x"08",
          2885 => x"55",
          2886 => x"89",
          2887 => x"75",
          2888 => x"d7",
          2889 => x"d8",
          2890 => x"9f",
          2891 => x"30",
          2892 => x"80",
          2893 => x"70",
          2894 => x"06",
          2895 => x"56",
          2896 => x"90",
          2897 => x"a4",
          2898 => x"98",
          2899 => x"78",
          2900 => x"3f",
          2901 => x"82",
          2902 => x"96",
          2903 => x"f7",
          2904 => x"02",
          2905 => x"05",
          2906 => x"ff",
          2907 => x"7c",
          2908 => x"fe",
          2909 => x"d6",
          2910 => x"cb",
          2911 => x"2e",
          2912 => x"81",
          2913 => x"bf",
          2914 => x"b8",
          2915 => x"b8",
          2916 => x"b8",
          2917 => x"c0",
          2918 => x"f2",
          2919 => x"82",
          2920 => x"52",
          2921 => x"51",
          2922 => x"3f",
          2923 => x"56",
          2924 => x"54",
          2925 => x"53",
          2926 => x"51",
          2927 => x"d6",
          2928 => x"83",
          2929 => x"78",
          2930 => x"0c",
          2931 => x"04",
          2932 => x"7f",
          2933 => x"8c",
          2934 => x"05",
          2935 => x"15",
          2936 => x"5c",
          2937 => x"5e",
          2938 => x"b6",
          2939 => x"b7",
          2940 => x"b6",
          2941 => x"b7",
          2942 => x"55",
          2943 => x"81",
          2944 => x"90",
          2945 => x"7b",
          2946 => x"38",
          2947 => x"74",
          2948 => x"7a",
          2949 => x"72",
          2950 => x"b6",
          2951 => x"b7",
          2952 => x"39",
          2953 => x"51",
          2954 => x"3f",
          2955 => x"80",
          2956 => x"18",
          2957 => x"27",
          2958 => x"08",
          2959 => x"e0",
          2960 => x"97",
          2961 => x"82",
          2962 => x"ff",
          2963 => x"84",
          2964 => x"39",
          2965 => x"72",
          2966 => x"38",
          2967 => x"82",
          2968 => x"ff",
          2969 => x"89",
          2970 => x"88",
          2971 => x"eb",
          2972 => x"55",
          2973 => x"08",
          2974 => x"d6",
          2975 => x"fc",
          2976 => x"8c",
          2977 => x"d3",
          2978 => x"74",
          2979 => x"c6",
          2980 => x"70",
          2981 => x"80",
          2982 => x"27",
          2983 => x"56",
          2984 => x"74",
          2985 => x"81",
          2986 => x"06",
          2987 => x"06",
          2988 => x"80",
          2989 => x"73",
          2990 => x"8a",
          2991 => x"bc",
          2992 => x"51",
          2993 => x"f2",
          2994 => x"a0",
          2995 => x"3f",
          2996 => x"ff",
          2997 => x"b7",
          2998 => x"8a",
          2999 => x"79",
          3000 => x"9c",
          3001 => x"d6",
          3002 => x"2b",
          3003 => x"51",
          3004 => x"2e",
          3005 => x"aa",
          3006 => x"3f",
          3007 => x"08",
          3008 => x"98",
          3009 => x"32",
          3010 => x"9b",
          3011 => x"70",
          3012 => x"75",
          3013 => x"58",
          3014 => x"51",
          3015 => x"24",
          3016 => x"9b",
          3017 => x"06",
          3018 => x"53",
          3019 => x"1e",
          3020 => x"26",
          3021 => x"ff",
          3022 => x"d6",
          3023 => x"3d",
          3024 => x"3d",
          3025 => x"05",
          3026 => x"94",
          3027 => x"98",
          3028 => x"b5",
          3029 => x"d4",
          3030 => x"a5",
          3031 => x"b7",
          3032 => x"b7",
          3033 => x"d4",
          3034 => x"82",
          3035 => x"ff",
          3036 => x"74",
          3037 => x"38",
          3038 => x"86",
          3039 => x"fe",
          3040 => x"c0",
          3041 => x"53",
          3042 => x"81",
          3043 => x"3f",
          3044 => x"51",
          3045 => x"80",
          3046 => x"3f",
          3047 => x"70",
          3048 => x"52",
          3049 => x"92",
          3050 => x"99",
          3051 => x"b7",
          3052 => x"b0",
          3053 => x"99",
          3054 => x"82",
          3055 => x"06",
          3056 => x"80",
          3057 => x"81",
          3058 => x"3f",
          3059 => x"51",
          3060 => x"80",
          3061 => x"3f",
          3062 => x"70",
          3063 => x"52",
          3064 => x"92",
          3065 => x"98",
          3066 => x"b8",
          3067 => x"f4",
          3068 => x"98",
          3069 => x"84",
          3070 => x"06",
          3071 => x"80",
          3072 => x"81",
          3073 => x"3f",
          3074 => x"51",
          3075 => x"80",
          3076 => x"3f",
          3077 => x"70",
          3078 => x"52",
          3079 => x"92",
          3080 => x"98",
          3081 => x"b8",
          3082 => x"b8",
          3083 => x"98",
          3084 => x"86",
          3085 => x"06",
          3086 => x"80",
          3087 => x"81",
          3088 => x"3f",
          3089 => x"51",
          3090 => x"80",
          3091 => x"3f",
          3092 => x"70",
          3093 => x"52",
          3094 => x"92",
          3095 => x"97",
          3096 => x"b8",
          3097 => x"fc",
          3098 => x"97",
          3099 => x"88",
          3100 => x"06",
          3101 => x"80",
          3102 => x"81",
          3103 => x"3f",
          3104 => x"51",
          3105 => x"80",
          3106 => x"3f",
          3107 => x"84",
          3108 => x"fb",
          3109 => x"02",
          3110 => x"05",
          3111 => x"56",
          3112 => x"75",
          3113 => x"3f",
          3114 => x"d0",
          3115 => x"73",
          3116 => x"53",
          3117 => x"52",
          3118 => x"51",
          3119 => x"3f",
          3120 => x"08",
          3121 => x"d6",
          3122 => x"80",
          3123 => x"31",
          3124 => x"73",
          3125 => x"d0",
          3126 => x"0b",
          3127 => x"33",
          3128 => x"2e",
          3129 => x"af",
          3130 => x"e8",
          3131 => x"75",
          3132 => x"c1",
          3133 => x"d8",
          3134 => x"8b",
          3135 => x"d8",
          3136 => x"e2",
          3137 => x"82",
          3138 => x"81",
          3139 => x"82",
          3140 => x"82",
          3141 => x"0b",
          3142 => x"c8",
          3143 => x"82",
          3144 => x"06",
          3145 => x"b9",
          3146 => x"52",
          3147 => x"d8",
          3148 => x"82",
          3149 => x"87",
          3150 => x"cd",
          3151 => x"70",
          3152 => x"7e",
          3153 => x"0c",
          3154 => x"7d",
          3155 => x"88",
          3156 => x"d8",
          3157 => x"06",
          3158 => x"2e",
          3159 => x"a3",
          3160 => x"59",
          3161 => x"b9",
          3162 => x"51",
          3163 => x"7d",
          3164 => x"82",
          3165 => x"81",
          3166 => x"82",
          3167 => x"7e",
          3168 => x"82",
          3169 => x"8d",
          3170 => x"70",
          3171 => x"ba",
          3172 => x"b0",
          3173 => x"3d",
          3174 => x"80",
          3175 => x"51",
          3176 => x"b5",
          3177 => x"05",
          3178 => x"3f",
          3179 => x"08",
          3180 => x"90",
          3181 => x"78",
          3182 => x"87",
          3183 => x"80",
          3184 => x"38",
          3185 => x"81",
          3186 => x"bd",
          3187 => x"78",
          3188 => x"ba",
          3189 => x"2e",
          3190 => x"8a",
          3191 => x"80",
          3192 => x"99",
          3193 => x"c0",
          3194 => x"38",
          3195 => x"82",
          3196 => x"bf",
          3197 => x"f9",
          3198 => x"38",
          3199 => x"24",
          3200 => x"80",
          3201 => x"8a",
          3202 => x"f8",
          3203 => x"38",
          3204 => x"78",
          3205 => x"8a",
          3206 => x"81",
          3207 => x"38",
          3208 => x"2e",
          3209 => x"8a",
          3210 => x"81",
          3211 => x"fd",
          3212 => x"39",
          3213 => x"80",
          3214 => x"84",
          3215 => x"ba",
          3216 => x"d8",
          3217 => x"fe",
          3218 => x"3d",
          3219 => x"53",
          3220 => x"51",
          3221 => x"82",
          3222 => x"80",
          3223 => x"38",
          3224 => x"f8",
          3225 => x"84",
          3226 => x"8e",
          3227 => x"d8",
          3228 => x"82",
          3229 => x"43",
          3230 => x"51",
          3231 => x"3f",
          3232 => x"5a",
          3233 => x"81",
          3234 => x"59",
          3235 => x"84",
          3236 => x"7a",
          3237 => x"38",
          3238 => x"b5",
          3239 => x"11",
          3240 => x"05",
          3241 => x"3f",
          3242 => x"08",
          3243 => x"de",
          3244 => x"fe",
          3245 => x"ff",
          3246 => x"eb",
          3247 => x"d6",
          3248 => x"2e",
          3249 => x"b5",
          3250 => x"11",
          3251 => x"05",
          3252 => x"3f",
          3253 => x"08",
          3254 => x"b2",
          3255 => x"94",
          3256 => x"f7",
          3257 => x"79",
          3258 => x"89",
          3259 => x"79",
          3260 => x"5b",
          3261 => x"62",
          3262 => x"eb",
          3263 => x"ff",
          3264 => x"ff",
          3265 => x"ea",
          3266 => x"d6",
          3267 => x"2e",
          3268 => x"b5",
          3269 => x"11",
          3270 => x"05",
          3271 => x"3f",
          3272 => x"08",
          3273 => x"e6",
          3274 => x"fe",
          3275 => x"ff",
          3276 => x"ea",
          3277 => x"d6",
          3278 => x"2e",
          3279 => x"82",
          3280 => x"ff",
          3281 => x"64",
          3282 => x"27",
          3283 => x"70",
          3284 => x"5e",
          3285 => x"7c",
          3286 => x"78",
          3287 => x"79",
          3288 => x"52",
          3289 => x"51",
          3290 => x"3f",
          3291 => x"81",
          3292 => x"d5",
          3293 => x"cc",
          3294 => x"92",
          3295 => x"ff",
          3296 => x"ff",
          3297 => x"e9",
          3298 => x"d6",
          3299 => x"df",
          3300 => x"b8",
          3301 => x"80",
          3302 => x"82",
          3303 => x"45",
          3304 => x"82",
          3305 => x"59",
          3306 => x"88",
          3307 => x"f8",
          3308 => x"39",
          3309 => x"33",
          3310 => x"2e",
          3311 => x"d4",
          3312 => x"ab",
          3313 => x"bb",
          3314 => x"80",
          3315 => x"82",
          3316 => x"45",
          3317 => x"d4",
          3318 => x"78",
          3319 => x"38",
          3320 => x"08",
          3321 => x"82",
          3322 => x"fc",
          3323 => x"b5",
          3324 => x"11",
          3325 => x"05",
          3326 => x"3f",
          3327 => x"08",
          3328 => x"82",
          3329 => x"59",
          3330 => x"89",
          3331 => x"f4",
          3332 => x"cc",
          3333 => x"b9",
          3334 => x"80",
          3335 => x"82",
          3336 => x"44",
          3337 => x"d4",
          3338 => x"78",
          3339 => x"38",
          3340 => x"08",
          3341 => x"82",
          3342 => x"59",
          3343 => x"88",
          3344 => x"8c",
          3345 => x"39",
          3346 => x"33",
          3347 => x"2e",
          3348 => x"d4",
          3349 => x"88",
          3350 => x"a0",
          3351 => x"44",
          3352 => x"f8",
          3353 => x"84",
          3354 => x"8e",
          3355 => x"d8",
          3356 => x"a7",
          3357 => x"5c",
          3358 => x"2e",
          3359 => x"5c",
          3360 => x"70",
          3361 => x"07",
          3362 => x"7f",
          3363 => x"5a",
          3364 => x"2e",
          3365 => x"a0",
          3366 => x"88",
          3367 => x"cc",
          3368 => x"3f",
          3369 => x"54",
          3370 => x"52",
          3371 => x"a0",
          3372 => x"d8",
          3373 => x"39",
          3374 => x"80",
          3375 => x"84",
          3376 => x"b6",
          3377 => x"d8",
          3378 => x"f9",
          3379 => x"3d",
          3380 => x"53",
          3381 => x"51",
          3382 => x"82",
          3383 => x"80",
          3384 => x"64",
          3385 => x"cf",
          3386 => x"34",
          3387 => x"45",
          3388 => x"fc",
          3389 => x"84",
          3390 => x"fe",
          3391 => x"d8",
          3392 => x"f9",
          3393 => x"70",
          3394 => x"82",
          3395 => x"ff",
          3396 => x"82",
          3397 => x"53",
          3398 => x"79",
          3399 => x"90",
          3400 => x"79",
          3401 => x"ae",
          3402 => x"38",
          3403 => x"9f",
          3404 => x"fe",
          3405 => x"ff",
          3406 => x"e6",
          3407 => x"d6",
          3408 => x"2e",
          3409 => x"59",
          3410 => x"05",
          3411 => x"64",
          3412 => x"ff",
          3413 => x"ba",
          3414 => x"8a",
          3415 => x"39",
          3416 => x"f4",
          3417 => x"84",
          3418 => x"bd",
          3419 => x"d8",
          3420 => x"f8",
          3421 => x"3d",
          3422 => x"53",
          3423 => x"51",
          3424 => x"82",
          3425 => x"80",
          3426 => x"61",
          3427 => x"c2",
          3428 => x"70",
          3429 => x"23",
          3430 => x"3d",
          3431 => x"53",
          3432 => x"51",
          3433 => x"82",
          3434 => x"df",
          3435 => x"39",
          3436 => x"54",
          3437 => x"f4",
          3438 => x"9f",
          3439 => x"b8",
          3440 => x"f8",
          3441 => x"ff",
          3442 => x"79",
          3443 => x"59",
          3444 => x"f7",
          3445 => x"9f",
          3446 => x"61",
          3447 => x"d0",
          3448 => x"fe",
          3449 => x"ff",
          3450 => x"df",
          3451 => x"d6",
          3452 => x"2e",
          3453 => x"59",
          3454 => x"05",
          3455 => x"82",
          3456 => x"78",
          3457 => x"39",
          3458 => x"51",
          3459 => x"ff",
          3460 => x"3d",
          3461 => x"53",
          3462 => x"51",
          3463 => x"82",
          3464 => x"80",
          3465 => x"38",
          3466 => x"f0",
          3467 => x"84",
          3468 => x"f5",
          3469 => x"d8",
          3470 => x"a0",
          3471 => x"71",
          3472 => x"84",
          3473 => x"3d",
          3474 => x"53",
          3475 => x"51",
          3476 => x"82",
          3477 => x"e5",
          3478 => x"39",
          3479 => x"54",
          3480 => x"80",
          3481 => x"f3",
          3482 => x"b8",
          3483 => x"f8",
          3484 => x"ff",
          3485 => x"79",
          3486 => x"59",
          3487 => x"f6",
          3488 => x"79",
          3489 => x"b5",
          3490 => x"11",
          3491 => x"05",
          3492 => x"3f",
          3493 => x"08",
          3494 => x"38",
          3495 => x"0c",
          3496 => x"05",
          3497 => x"39",
          3498 => x"51",
          3499 => x"ff",
          3500 => x"3d",
          3501 => x"53",
          3502 => x"51",
          3503 => x"82",
          3504 => x"80",
          3505 => x"38",
          3506 => x"bb",
          3507 => x"a6",
          3508 => x"59",
          3509 => x"3d",
          3510 => x"53",
          3511 => x"51",
          3512 => x"82",
          3513 => x"80",
          3514 => x"38",
          3515 => x"bb",
          3516 => x"a5",
          3517 => x"59",
          3518 => x"d6",
          3519 => x"2e",
          3520 => x"82",
          3521 => x"52",
          3522 => x"51",
          3523 => x"3f",
          3524 => x"82",
          3525 => x"c1",
          3526 => x"a5",
          3527 => x"ee",
          3528 => x"80",
          3529 => x"3f",
          3530 => x"a8",
          3531 => x"3f",
          3532 => x"97",
          3533 => x"78",
          3534 => x"d2",
          3535 => x"52",
          3536 => x"f8",
          3537 => x"d8",
          3538 => x"d6",
          3539 => x"2e",
          3540 => x"82",
          3541 => x"46",
          3542 => x"84",
          3543 => x"e5",
          3544 => x"d8",
          3545 => x"06",
          3546 => x"80",
          3547 => x"38",
          3548 => x"08",
          3549 => x"3f",
          3550 => x"08",
          3551 => x"c1",
          3552 => x"7a",
          3553 => x"38",
          3554 => x"89",
          3555 => x"2e",
          3556 => x"ca",
          3557 => x"2e",
          3558 => x"c2",
          3559 => x"94",
          3560 => x"82",
          3561 => x"80",
          3562 => x"9c",
          3563 => x"ff",
          3564 => x"ff",
          3565 => x"b8",
          3566 => x"b5",
          3567 => x"05",
          3568 => x"3f",
          3569 => x"55",
          3570 => x"54",
          3571 => x"bc",
          3572 => x"3d",
          3573 => x"51",
          3574 => x"3f",
          3575 => x"54",
          3576 => x"bc",
          3577 => x"3d",
          3578 => x"51",
          3579 => x"3f",
          3580 => x"58",
          3581 => x"57",
          3582 => x"55",
          3583 => x"80",
          3584 => x"80",
          3585 => x"3d",
          3586 => x"51",
          3587 => x"82",
          3588 => x"82",
          3589 => x"09",
          3590 => x"72",
          3591 => x"51",
          3592 => x"80",
          3593 => x"26",
          3594 => x"5a",
          3595 => x"59",
          3596 => x"8d",
          3597 => x"70",
          3598 => x"5c",
          3599 => x"c3",
          3600 => x"32",
          3601 => x"07",
          3602 => x"38",
          3603 => x"09",
          3604 => x"38",
          3605 => x"51",
          3606 => x"3f",
          3607 => x"f5",
          3608 => x"39",
          3609 => x"51",
          3610 => x"3f",
          3611 => x"f6",
          3612 => x"0b",
          3613 => x"34",
          3614 => x"8c",
          3615 => x"84",
          3616 => x"51",
          3617 => x"82",
          3618 => x"90",
          3619 => x"94",
          3620 => x"53",
          3621 => x"52",
          3622 => x"95",
          3623 => x"d6",
          3624 => x"87",
          3625 => x"0c",
          3626 => x"9c",
          3627 => x"84",
          3628 => x"51",
          3629 => x"82",
          3630 => x"90",
          3631 => x"94",
          3632 => x"53",
          3633 => x"52",
          3634 => x"e5",
          3635 => x"d6",
          3636 => x"87",
          3637 => x"0c",
          3638 => x"0b",
          3639 => x"84",
          3640 => x"83",
          3641 => x"94",
          3642 => x"a0",
          3643 => x"80",
          3644 => x"05",
          3645 => x"a0",
          3646 => x"27",
          3647 => x"a0",
          3648 => x"87",
          3649 => x"f1",
          3650 => x"05",
          3651 => x"a0",
          3652 => x"27",
          3653 => x"52",
          3654 => x"a7",
          3655 => x"52",
          3656 => x"a7",
          3657 => x"52",
          3658 => x"a7",
          3659 => x"52",
          3660 => x"a7",
          3661 => x"52",
          3662 => x"a6",
          3663 => x"52",
          3664 => x"f7",
          3665 => x"be",
          3666 => x"3f",
          3667 => x"59",
          3668 => x"5a",
          3669 => x"05",
          3670 => x"80",
          3671 => x"70",
          3672 => x"0c",
          3673 => x"b8",
          3674 => x"bc",
          3675 => x"fc",
          3676 => x"f2",
          3677 => x"3f",
          3678 => x"82",
          3679 => x"ff",
          3680 => x"82",
          3681 => x"ff",
          3682 => x"80",
          3683 => x"91",
          3684 => x"51",
          3685 => x"ef",
          3686 => x"04",
          3687 => x"80",
          3688 => x"71",
          3689 => x"86",
          3690 => x"d6",
          3691 => x"ff",
          3692 => x"ff",
          3693 => x"72",
          3694 => x"38",
          3695 => x"d8",
          3696 => x"0d",
          3697 => x"0d",
          3698 => x"54",
          3699 => x"52",
          3700 => x"2e",
          3701 => x"72",
          3702 => x"a0",
          3703 => x"06",
          3704 => x"13",
          3705 => x"72",
          3706 => x"a2",
          3707 => x"06",
          3708 => x"13",
          3709 => x"72",
          3710 => x"2e",
          3711 => x"9f",
          3712 => x"81",
          3713 => x"72",
          3714 => x"70",
          3715 => x"38",
          3716 => x"80",
          3717 => x"73",
          3718 => x"39",
          3719 => x"80",
          3720 => x"54",
          3721 => x"83",
          3722 => x"70",
          3723 => x"38",
          3724 => x"80",
          3725 => x"54",
          3726 => x"09",
          3727 => x"38",
          3728 => x"a2",
          3729 => x"70",
          3730 => x"07",
          3731 => x"70",
          3732 => x"38",
          3733 => x"81",
          3734 => x"71",
          3735 => x"51",
          3736 => x"d8",
          3737 => x"0d",
          3738 => x"0d",
          3739 => x"08",
          3740 => x"38",
          3741 => x"05",
          3742 => x"d6",
          3743 => x"d6",
          3744 => x"38",
          3745 => x"39",
          3746 => x"82",
          3747 => x"86",
          3748 => x"fc",
          3749 => x"82",
          3750 => x"05",
          3751 => x"52",
          3752 => x"81",
          3753 => x"13",
          3754 => x"51",
          3755 => x"9e",
          3756 => x"38",
          3757 => x"51",
          3758 => x"97",
          3759 => x"38",
          3760 => x"51",
          3761 => x"bb",
          3762 => x"38",
          3763 => x"51",
          3764 => x"bb",
          3765 => x"38",
          3766 => x"55",
          3767 => x"87",
          3768 => x"d9",
          3769 => x"22",
          3770 => x"73",
          3771 => x"80",
          3772 => x"0b",
          3773 => x"9c",
          3774 => x"87",
          3775 => x"0c",
          3776 => x"87",
          3777 => x"0c",
          3778 => x"87",
          3779 => x"0c",
          3780 => x"87",
          3781 => x"0c",
          3782 => x"87",
          3783 => x"0c",
          3784 => x"87",
          3785 => x"0c",
          3786 => x"98",
          3787 => x"87",
          3788 => x"0c",
          3789 => x"c0",
          3790 => x"80",
          3791 => x"d6",
          3792 => x"3d",
          3793 => x"3d",
          3794 => x"87",
          3795 => x"5d",
          3796 => x"87",
          3797 => x"08",
          3798 => x"23",
          3799 => x"b8",
          3800 => x"82",
          3801 => x"c0",
          3802 => x"5a",
          3803 => x"34",
          3804 => x"b0",
          3805 => x"84",
          3806 => x"c0",
          3807 => x"5a",
          3808 => x"34",
          3809 => x"a8",
          3810 => x"86",
          3811 => x"c0",
          3812 => x"5c",
          3813 => x"23",
          3814 => x"a0",
          3815 => x"8a",
          3816 => x"7d",
          3817 => x"ff",
          3818 => x"7b",
          3819 => x"06",
          3820 => x"33",
          3821 => x"33",
          3822 => x"33",
          3823 => x"33",
          3824 => x"33",
          3825 => x"ff",
          3826 => x"82",
          3827 => x"ff",
          3828 => x"8f",
          3829 => x"fb",
          3830 => x"9f",
          3831 => x"d3",
          3832 => x"81",
          3833 => x"55",
          3834 => x"94",
          3835 => x"80",
          3836 => x"87",
          3837 => x"51",
          3838 => x"96",
          3839 => x"06",
          3840 => x"70",
          3841 => x"38",
          3842 => x"70",
          3843 => x"51",
          3844 => x"72",
          3845 => x"81",
          3846 => x"70",
          3847 => x"38",
          3848 => x"70",
          3849 => x"51",
          3850 => x"38",
          3851 => x"06",
          3852 => x"94",
          3853 => x"80",
          3854 => x"87",
          3855 => x"52",
          3856 => x"74",
          3857 => x"0c",
          3858 => x"04",
          3859 => x"02",
          3860 => x"70",
          3861 => x"2a",
          3862 => x"70",
          3863 => x"34",
          3864 => x"04",
          3865 => x"79",
          3866 => x"33",
          3867 => x"06",
          3868 => x"70",
          3869 => x"fc",
          3870 => x"ff",
          3871 => x"82",
          3872 => x"70",
          3873 => x"59",
          3874 => x"87",
          3875 => x"51",
          3876 => x"86",
          3877 => x"94",
          3878 => x"08",
          3879 => x"70",
          3880 => x"54",
          3881 => x"2e",
          3882 => x"91",
          3883 => x"06",
          3884 => x"d7",
          3885 => x"32",
          3886 => x"51",
          3887 => x"2e",
          3888 => x"93",
          3889 => x"06",
          3890 => x"ff",
          3891 => x"81",
          3892 => x"87",
          3893 => x"52",
          3894 => x"86",
          3895 => x"94",
          3896 => x"72",
          3897 => x"74",
          3898 => x"ff",
          3899 => x"57",
          3900 => x"38",
          3901 => x"d8",
          3902 => x"0d",
          3903 => x"0d",
          3904 => x"33",
          3905 => x"06",
          3906 => x"c0",
          3907 => x"72",
          3908 => x"38",
          3909 => x"94",
          3910 => x"70",
          3911 => x"81",
          3912 => x"51",
          3913 => x"e2",
          3914 => x"ff",
          3915 => x"c0",
          3916 => x"70",
          3917 => x"38",
          3918 => x"90",
          3919 => x"70",
          3920 => x"82",
          3921 => x"51",
          3922 => x"04",
          3923 => x"82",
          3924 => x"70",
          3925 => x"52",
          3926 => x"94",
          3927 => x"80",
          3928 => x"87",
          3929 => x"52",
          3930 => x"82",
          3931 => x"06",
          3932 => x"ff",
          3933 => x"2e",
          3934 => x"81",
          3935 => x"87",
          3936 => x"52",
          3937 => x"86",
          3938 => x"94",
          3939 => x"08",
          3940 => x"70",
          3941 => x"53",
          3942 => x"d6",
          3943 => x"3d",
          3944 => x"3d",
          3945 => x"9e",
          3946 => x"9c",
          3947 => x"51",
          3948 => x"2e",
          3949 => x"87",
          3950 => x"08",
          3951 => x"0c",
          3952 => x"a8",
          3953 => x"f4",
          3954 => x"9e",
          3955 => x"d3",
          3956 => x"c0",
          3957 => x"82",
          3958 => x"87",
          3959 => x"08",
          3960 => x"0c",
          3961 => x"a0",
          3962 => x"84",
          3963 => x"9e",
          3964 => x"d4",
          3965 => x"c0",
          3966 => x"82",
          3967 => x"87",
          3968 => x"08",
          3969 => x"0c",
          3970 => x"b8",
          3971 => x"94",
          3972 => x"9e",
          3973 => x"d4",
          3974 => x"c0",
          3975 => x"82",
          3976 => x"87",
          3977 => x"08",
          3978 => x"0c",
          3979 => x"80",
          3980 => x"82",
          3981 => x"87",
          3982 => x"08",
          3983 => x"0c",
          3984 => x"88",
          3985 => x"ac",
          3986 => x"9e",
          3987 => x"d4",
          3988 => x"0b",
          3989 => x"34",
          3990 => x"c0",
          3991 => x"70",
          3992 => x"06",
          3993 => x"70",
          3994 => x"38",
          3995 => x"82",
          3996 => x"80",
          3997 => x"9e",
          3998 => x"88",
          3999 => x"51",
          4000 => x"80",
          4001 => x"81",
          4002 => x"d4",
          4003 => x"0b",
          4004 => x"90",
          4005 => x"80",
          4006 => x"52",
          4007 => x"2e",
          4008 => x"52",
          4009 => x"b7",
          4010 => x"87",
          4011 => x"08",
          4012 => x"80",
          4013 => x"52",
          4014 => x"83",
          4015 => x"71",
          4016 => x"34",
          4017 => x"c0",
          4018 => x"70",
          4019 => x"06",
          4020 => x"70",
          4021 => x"38",
          4022 => x"82",
          4023 => x"80",
          4024 => x"9e",
          4025 => x"90",
          4026 => x"51",
          4027 => x"80",
          4028 => x"81",
          4029 => x"d4",
          4030 => x"0b",
          4031 => x"90",
          4032 => x"80",
          4033 => x"52",
          4034 => x"2e",
          4035 => x"52",
          4036 => x"bb",
          4037 => x"87",
          4038 => x"08",
          4039 => x"80",
          4040 => x"52",
          4041 => x"83",
          4042 => x"71",
          4043 => x"34",
          4044 => x"c0",
          4045 => x"70",
          4046 => x"06",
          4047 => x"70",
          4048 => x"38",
          4049 => x"82",
          4050 => x"80",
          4051 => x"9e",
          4052 => x"80",
          4053 => x"51",
          4054 => x"80",
          4055 => x"81",
          4056 => x"d4",
          4057 => x"0b",
          4058 => x"90",
          4059 => x"80",
          4060 => x"52",
          4061 => x"83",
          4062 => x"71",
          4063 => x"34",
          4064 => x"90",
          4065 => x"80",
          4066 => x"2a",
          4067 => x"70",
          4068 => x"34",
          4069 => x"c0",
          4070 => x"70",
          4071 => x"51",
          4072 => x"80",
          4073 => x"81",
          4074 => x"d4",
          4075 => x"c0",
          4076 => x"70",
          4077 => x"70",
          4078 => x"51",
          4079 => x"d4",
          4080 => x"0b",
          4081 => x"90",
          4082 => x"06",
          4083 => x"70",
          4084 => x"38",
          4085 => x"82",
          4086 => x"87",
          4087 => x"08",
          4088 => x"51",
          4089 => x"d4",
          4090 => x"3d",
          4091 => x"3d",
          4092 => x"c8",
          4093 => x"e3",
          4094 => x"b4",
          4095 => x"80",
          4096 => x"82",
          4097 => x"ff",
          4098 => x"82",
          4099 => x"ff",
          4100 => x"82",
          4101 => x"54",
          4102 => x"94",
          4103 => x"90",
          4104 => x"94",
          4105 => x"52",
          4106 => x"51",
          4107 => x"3f",
          4108 => x"33",
          4109 => x"2e",
          4110 => x"d4",
          4111 => x"d4",
          4112 => x"54",
          4113 => x"a4",
          4114 => x"8f",
          4115 => x"b8",
          4116 => x"80",
          4117 => x"82",
          4118 => x"82",
          4119 => x"11",
          4120 => x"be",
          4121 => x"92",
          4122 => x"d4",
          4123 => x"73",
          4124 => x"38",
          4125 => x"08",
          4126 => x"08",
          4127 => x"82",
          4128 => x"ff",
          4129 => x"82",
          4130 => x"54",
          4131 => x"94",
          4132 => x"80",
          4133 => x"84",
          4134 => x"52",
          4135 => x"51",
          4136 => x"3f",
          4137 => x"33",
          4138 => x"2e",
          4139 => x"d4",
          4140 => x"82",
          4141 => x"ff",
          4142 => x"82",
          4143 => x"54",
          4144 => x"8e",
          4145 => x"c4",
          4146 => x"bf",
          4147 => x"92",
          4148 => x"d4",
          4149 => x"73",
          4150 => x"38",
          4151 => x"33",
          4152 => x"d4",
          4153 => x"f3",
          4154 => x"b5",
          4155 => x"80",
          4156 => x"82",
          4157 => x"ff",
          4158 => x"82",
          4159 => x"54",
          4160 => x"89",
          4161 => x"88",
          4162 => x"da",
          4163 => x"bc",
          4164 => x"80",
          4165 => x"82",
          4166 => x"ff",
          4167 => x"82",
          4168 => x"54",
          4169 => x"89",
          4170 => x"a0",
          4171 => x"b6",
          4172 => x"be",
          4173 => x"80",
          4174 => x"82",
          4175 => x"ff",
          4176 => x"82",
          4177 => x"ff",
          4178 => x"82",
          4179 => x"52",
          4180 => x"51",
          4181 => x"3f",
          4182 => x"08",
          4183 => x"e4",
          4184 => x"f7",
          4185 => x"a0",
          4186 => x"c1",
          4187 => x"90",
          4188 => x"c1",
          4189 => x"ac",
          4190 => x"d4",
          4191 => x"82",
          4192 => x"ff",
          4193 => x"82",
          4194 => x"56",
          4195 => x"52",
          4196 => x"9d",
          4197 => x"d8",
          4198 => x"c0",
          4199 => x"31",
          4200 => x"d6",
          4201 => x"82",
          4202 => x"ff",
          4203 => x"82",
          4204 => x"54",
          4205 => x"a9",
          4206 => x"ac",
          4207 => x"84",
          4208 => x"51",
          4209 => x"82",
          4210 => x"bd",
          4211 => x"76",
          4212 => x"54",
          4213 => x"08",
          4214 => x"90",
          4215 => x"fb",
          4216 => x"b6",
          4217 => x"80",
          4218 => x"82",
          4219 => x"56",
          4220 => x"52",
          4221 => x"b9",
          4222 => x"d8",
          4223 => x"c0",
          4224 => x"31",
          4225 => x"d6",
          4226 => x"82",
          4227 => x"ff",
          4228 => x"8a",
          4229 => x"f0",
          4230 => x"0d",
          4231 => x"0d",
          4232 => x"33",
          4233 => x"71",
          4234 => x"38",
          4235 => x"82",
          4236 => x"52",
          4237 => x"82",
          4238 => x"9d",
          4239 => x"f0",
          4240 => x"82",
          4241 => x"91",
          4242 => x"80",
          4243 => x"82",
          4244 => x"85",
          4245 => x"8c",
          4246 => x"ff",
          4247 => x"0d",
          4248 => x"80",
          4249 => x"0b",
          4250 => x"84",
          4251 => x"d4",
          4252 => x"c0",
          4253 => x"04",
          4254 => x"76",
          4255 => x"98",
          4256 => x"2b",
          4257 => x"72",
          4258 => x"82",
          4259 => x"51",
          4260 => x"80",
          4261 => x"98",
          4262 => x"53",
          4263 => x"9c",
          4264 => x"94",
          4265 => x"02",
          4266 => x"05",
          4267 => x"52",
          4268 => x"72",
          4269 => x"06",
          4270 => x"53",
          4271 => x"d8",
          4272 => x"0d",
          4273 => x"0d",
          4274 => x"05",
          4275 => x"71",
          4276 => x"54",
          4277 => x"b1",
          4278 => x"bc",
          4279 => x"51",
          4280 => x"3f",
          4281 => x"08",
          4282 => x"ff",
          4283 => x"82",
          4284 => x"52",
          4285 => x"ad",
          4286 => x"33",
          4287 => x"72",
          4288 => x"81",
          4289 => x"cc",
          4290 => x"ff",
          4291 => x"74",
          4292 => x"3d",
          4293 => x"3d",
          4294 => x"84",
          4295 => x"33",
          4296 => x"bb",
          4297 => x"d5",
          4298 => x"84",
          4299 => x"cc",
          4300 => x"51",
          4301 => x"58",
          4302 => x"2e",
          4303 => x"51",
          4304 => x"82",
          4305 => x"70",
          4306 => x"d4",
          4307 => x"19",
          4308 => x"56",
          4309 => x"3f",
          4310 => x"08",
          4311 => x"d5",
          4312 => x"84",
          4313 => x"cc",
          4314 => x"51",
          4315 => x"80",
          4316 => x"75",
          4317 => x"74",
          4318 => x"ec",
          4319 => x"a4",
          4320 => x"55",
          4321 => x"a4",
          4322 => x"ff",
          4323 => x"75",
          4324 => x"80",
          4325 => x"a4",
          4326 => x"2e",
          4327 => x"d5",
          4328 => x"75",
          4329 => x"38",
          4330 => x"33",
          4331 => x"38",
          4332 => x"05",
          4333 => x"78",
          4334 => x"80",
          4335 => x"82",
          4336 => x"52",
          4337 => x"a2",
          4338 => x"d5",
          4339 => x"80",
          4340 => x"8c",
          4341 => x"fd",
          4342 => x"d4",
          4343 => x"54",
          4344 => x"71",
          4345 => x"38",
          4346 => x"e9",
          4347 => x"0c",
          4348 => x"14",
          4349 => x"80",
          4350 => x"80",
          4351 => x"a4",
          4352 => x"a0",
          4353 => x"80",
          4354 => x"71",
          4355 => x"9f",
          4356 => x"a0",
          4357 => x"bd",
          4358 => x"82",
          4359 => x"85",
          4360 => x"dc",
          4361 => x"57",
          4362 => x"d5",
          4363 => x"80",
          4364 => x"82",
          4365 => x"80",
          4366 => x"d5",
          4367 => x"80",
          4368 => x"3d",
          4369 => x"81",
          4370 => x"82",
          4371 => x"80",
          4372 => x"75",
          4373 => x"b0",
          4374 => x"d8",
          4375 => x"0b",
          4376 => x"08",
          4377 => x"82",
          4378 => x"ff",
          4379 => x"55",
          4380 => x"34",
          4381 => x"52",
          4382 => x"c6",
          4383 => x"ff",
          4384 => x"74",
          4385 => x"81",
          4386 => x"38",
          4387 => x"04",
          4388 => x"aa",
          4389 => x"3d",
          4390 => x"81",
          4391 => x"80",
          4392 => x"a0",
          4393 => x"f5",
          4394 => x"d6",
          4395 => x"95",
          4396 => x"82",
          4397 => x"54",
          4398 => x"52",
          4399 => x"52",
          4400 => x"f1",
          4401 => x"d8",
          4402 => x"a5",
          4403 => x"ff",
          4404 => x"82",
          4405 => x"81",
          4406 => x"80",
          4407 => x"d8",
          4408 => x"38",
          4409 => x"08",
          4410 => x"17",
          4411 => x"74",
          4412 => x"70",
          4413 => x"07",
          4414 => x"55",
          4415 => x"2e",
          4416 => x"ff",
          4417 => x"d5",
          4418 => x"11",
          4419 => x"80",
          4420 => x"82",
          4421 => x"80",
          4422 => x"82",
          4423 => x"ff",
          4424 => x"78",
          4425 => x"81",
          4426 => x"75",
          4427 => x"ff",
          4428 => x"79",
          4429 => x"d0",
          4430 => x"08",
          4431 => x"d8",
          4432 => x"80",
          4433 => x"d6",
          4434 => x"3d",
          4435 => x"3d",
          4436 => x"71",
          4437 => x"33",
          4438 => x"58",
          4439 => x"09",
          4440 => x"38",
          4441 => x"05",
          4442 => x"27",
          4443 => x"17",
          4444 => x"71",
          4445 => x"55",
          4446 => x"09",
          4447 => x"38",
          4448 => x"ea",
          4449 => x"73",
          4450 => x"d5",
          4451 => x"08",
          4452 => x"b0",
          4453 => x"d6",
          4454 => x"79",
          4455 => x"51",
          4456 => x"3f",
          4457 => x"08",
          4458 => x"84",
          4459 => x"74",
          4460 => x"38",
          4461 => x"88",
          4462 => x"fc",
          4463 => x"39",
          4464 => x"8c",
          4465 => x"53",
          4466 => x"c5",
          4467 => x"d6",
          4468 => x"2e",
          4469 => x"1b",
          4470 => x"77",
          4471 => x"3f",
          4472 => x"08",
          4473 => x"55",
          4474 => x"74",
          4475 => x"81",
          4476 => x"ff",
          4477 => x"82",
          4478 => x"8b",
          4479 => x"73",
          4480 => x"0c",
          4481 => x"04",
          4482 => x"b0",
          4483 => x"3d",
          4484 => x"08",
          4485 => x"80",
          4486 => x"34",
          4487 => x"33",
          4488 => x"08",
          4489 => x"81",
          4490 => x"82",
          4491 => x"55",
          4492 => x"38",
          4493 => x"80",
          4494 => x"38",
          4495 => x"06",
          4496 => x"80",
          4497 => x"38",
          4498 => x"9f",
          4499 => x"d8",
          4500 => x"a0",
          4501 => x"d8",
          4502 => x"81",
          4503 => x"53",
          4504 => x"d6",
          4505 => x"80",
          4506 => x"82",
          4507 => x"80",
          4508 => x"82",
          4509 => x"ff",
          4510 => x"80",
          4511 => x"d6",
          4512 => x"82",
          4513 => x"53",
          4514 => x"90",
          4515 => x"54",
          4516 => x"3f",
          4517 => x"08",
          4518 => x"d8",
          4519 => x"09",
          4520 => x"d0",
          4521 => x"d8",
          4522 => x"ae",
          4523 => x"d6",
          4524 => x"80",
          4525 => x"d8",
          4526 => x"38",
          4527 => x"08",
          4528 => x"17",
          4529 => x"74",
          4530 => x"74",
          4531 => x"52",
          4532 => x"c2",
          4533 => x"70",
          4534 => x"5c",
          4535 => x"27",
          4536 => x"5b",
          4537 => x"09",
          4538 => x"97",
          4539 => x"75",
          4540 => x"34",
          4541 => x"82",
          4542 => x"80",
          4543 => x"f9",
          4544 => x"3d",
          4545 => x"3f",
          4546 => x"08",
          4547 => x"98",
          4548 => x"78",
          4549 => x"38",
          4550 => x"06",
          4551 => x"33",
          4552 => x"70",
          4553 => x"ee",
          4554 => x"98",
          4555 => x"2c",
          4556 => x"05",
          4557 => x"82",
          4558 => x"70",
          4559 => x"33",
          4560 => x"51",
          4561 => x"59",
          4562 => x"56",
          4563 => x"80",
          4564 => x"74",
          4565 => x"74",
          4566 => x"29",
          4567 => x"05",
          4568 => x"51",
          4569 => x"24",
          4570 => x"76",
          4571 => x"77",
          4572 => x"3f",
          4573 => x"08",
          4574 => x"54",
          4575 => x"d7",
          4576 => x"ee",
          4577 => x"56",
          4578 => x"81",
          4579 => x"81",
          4580 => x"70",
          4581 => x"81",
          4582 => x"51",
          4583 => x"26",
          4584 => x"53",
          4585 => x"51",
          4586 => x"82",
          4587 => x"81",
          4588 => x"73",
          4589 => x"39",
          4590 => x"80",
          4591 => x"38",
          4592 => x"74",
          4593 => x"34",
          4594 => x"70",
          4595 => x"ee",
          4596 => x"98",
          4597 => x"2c",
          4598 => x"70",
          4599 => x"c3",
          4600 => x"5e",
          4601 => x"57",
          4602 => x"74",
          4603 => x"81",
          4604 => x"38",
          4605 => x"14",
          4606 => x"80",
          4607 => x"94",
          4608 => x"82",
          4609 => x"92",
          4610 => x"ee",
          4611 => x"82",
          4612 => x"78",
          4613 => x"75",
          4614 => x"54",
          4615 => x"fd",
          4616 => x"84",
          4617 => x"c0",
          4618 => x"08",
          4619 => x"9c",
          4620 => x"7e",
          4621 => x"38",
          4622 => x"33",
          4623 => x"27",
          4624 => x"98",
          4625 => x"2c",
          4626 => x"75",
          4627 => x"74",
          4628 => x"33",
          4629 => x"74",
          4630 => x"29",
          4631 => x"05",
          4632 => x"82",
          4633 => x"56",
          4634 => x"39",
          4635 => x"33",
          4636 => x"54",
          4637 => x"9c",
          4638 => x"54",
          4639 => x"74",
          4640 => x"98",
          4641 => x"7e",
          4642 => x"81",
          4643 => x"82",
          4644 => x"82",
          4645 => x"70",
          4646 => x"29",
          4647 => x"05",
          4648 => x"82",
          4649 => x"5a",
          4650 => x"74",
          4651 => x"38",
          4652 => x"08",
          4653 => x"70",
          4654 => x"ff",
          4655 => x"74",
          4656 => x"29",
          4657 => x"05",
          4658 => x"82",
          4659 => x"56",
          4660 => x"75",
          4661 => x"82",
          4662 => x"70",
          4663 => x"98",
          4664 => x"98",
          4665 => x"56",
          4666 => x"25",
          4667 => x"82",
          4668 => x"52",
          4669 => x"a1",
          4670 => x"81",
          4671 => x"81",
          4672 => x"70",
          4673 => x"ee",
          4674 => x"51",
          4675 => x"24",
          4676 => x"ee",
          4677 => x"34",
          4678 => x"1b",
          4679 => x"9c",
          4680 => x"82",
          4681 => x"f3",
          4682 => x"fd",
          4683 => x"9c",
          4684 => x"ff",
          4685 => x"73",
          4686 => x"c6",
          4687 => x"98",
          4688 => x"54",
          4689 => x"98",
          4690 => x"54",
          4691 => x"9c",
          4692 => x"bc",
          4693 => x"51",
          4694 => x"3f",
          4695 => x"33",
          4696 => x"70",
          4697 => x"ee",
          4698 => x"51",
          4699 => x"74",
          4700 => x"74",
          4701 => x"14",
          4702 => x"82",
          4703 => x"52",
          4704 => x"ff",
          4705 => x"74",
          4706 => x"29",
          4707 => x"05",
          4708 => x"82",
          4709 => x"58",
          4710 => x"75",
          4711 => x"82",
          4712 => x"52",
          4713 => x"a0",
          4714 => x"ee",
          4715 => x"98",
          4716 => x"2c",
          4717 => x"33",
          4718 => x"57",
          4719 => x"fa",
          4720 => x"f2",
          4721 => x"88",
          4722 => x"e9",
          4723 => x"80",
          4724 => x"80",
          4725 => x"98",
          4726 => x"98",
          4727 => x"55",
          4728 => x"de",
          4729 => x"39",
          4730 => x"33",
          4731 => x"80",
          4732 => x"f2",
          4733 => x"8a",
          4734 => x"b9",
          4735 => x"98",
          4736 => x"f6",
          4737 => x"d6",
          4738 => x"ff",
          4739 => x"96",
          4740 => x"98",
          4741 => x"80",
          4742 => x"81",
          4743 => x"79",
          4744 => x"3f",
          4745 => x"7a",
          4746 => x"82",
          4747 => x"80",
          4748 => x"98",
          4749 => x"d6",
          4750 => x"3d",
          4751 => x"ee",
          4752 => x"73",
          4753 => x"ba",
          4754 => x"bc",
          4755 => x"51",
          4756 => x"3f",
          4757 => x"33",
          4758 => x"73",
          4759 => x"34",
          4760 => x"06",
          4761 => x"82",
          4762 => x"82",
          4763 => x"55",
          4764 => x"2e",
          4765 => x"ff",
          4766 => x"82",
          4767 => x"74",
          4768 => x"98",
          4769 => x"ff",
          4770 => x"55",
          4771 => x"ad",
          4772 => x"54",
          4773 => x"74",
          4774 => x"bc",
          4775 => x"33",
          4776 => x"91",
          4777 => x"80",
          4778 => x"80",
          4779 => x"98",
          4780 => x"98",
          4781 => x"55",
          4782 => x"d5",
          4783 => x"bc",
          4784 => x"51",
          4785 => x"3f",
          4786 => x"33",
          4787 => x"70",
          4788 => x"ee",
          4789 => x"51",
          4790 => x"74",
          4791 => x"38",
          4792 => x"08",
          4793 => x"ff",
          4794 => x"74",
          4795 => x"29",
          4796 => x"05",
          4797 => x"82",
          4798 => x"58",
          4799 => x"75",
          4800 => x"f7",
          4801 => x"ee",
          4802 => x"81",
          4803 => x"ee",
          4804 => x"56",
          4805 => x"27",
          4806 => x"82",
          4807 => x"52",
          4808 => x"73",
          4809 => x"34",
          4810 => x"33",
          4811 => x"9d",
          4812 => x"ee",
          4813 => x"81",
          4814 => x"ee",
          4815 => x"56",
          4816 => x"26",
          4817 => x"ba",
          4818 => x"9c",
          4819 => x"82",
          4820 => x"ee",
          4821 => x"0b",
          4822 => x"34",
          4823 => x"ee",
          4824 => x"9e",
          4825 => x"38",
          4826 => x"08",
          4827 => x"2e",
          4828 => x"51",
          4829 => x"3f",
          4830 => x"08",
          4831 => x"34",
          4832 => x"08",
          4833 => x"81",
          4834 => x"52",
          4835 => x"a6",
          4836 => x"5b",
          4837 => x"7a",
          4838 => x"d4",
          4839 => x"11",
          4840 => x"74",
          4841 => x"38",
          4842 => x"a4",
          4843 => x"d6",
          4844 => x"ee",
          4845 => x"d6",
          4846 => x"ff",
          4847 => x"53",
          4848 => x"51",
          4849 => x"3f",
          4850 => x"80",
          4851 => x"08",
          4852 => x"2e",
          4853 => x"74",
          4854 => x"ac",
          4855 => x"7a",
          4856 => x"81",
          4857 => x"82",
          4858 => x"55",
          4859 => x"a4",
          4860 => x"ff",
          4861 => x"82",
          4862 => x"82",
          4863 => x"82",
          4864 => x"81",
          4865 => x"05",
          4866 => x"79",
          4867 => x"d8",
          4868 => x"39",
          4869 => x"82",
          4870 => x"70",
          4871 => x"74",
          4872 => x"38",
          4873 => x"a3",
          4874 => x"d6",
          4875 => x"ee",
          4876 => x"d6",
          4877 => x"ff",
          4878 => x"53",
          4879 => x"51",
          4880 => x"3f",
          4881 => x"73",
          4882 => x"5b",
          4883 => x"82",
          4884 => x"74",
          4885 => x"ee",
          4886 => x"ee",
          4887 => x"79",
          4888 => x"3f",
          4889 => x"82",
          4890 => x"70",
          4891 => x"82",
          4892 => x"59",
          4893 => x"77",
          4894 => x"38",
          4895 => x"08",
          4896 => x"54",
          4897 => x"9c",
          4898 => x"70",
          4899 => x"ff",
          4900 => x"f4",
          4901 => x"ee",
          4902 => x"73",
          4903 => x"e2",
          4904 => x"bc",
          4905 => x"51",
          4906 => x"3f",
          4907 => x"33",
          4908 => x"73",
          4909 => x"34",
          4910 => x"ff",
          4911 => x"8f",
          4912 => x"71",
          4913 => x"81",
          4914 => x"82",
          4915 => x"81",
          4916 => x"c4",
          4917 => x"82",
          4918 => x"25",
          4919 => x"0b",
          4920 => x"0c",
          4921 => x"d6",
          4922 => x"d6",
          4923 => x"29",
          4924 => x"08",
          4925 => x"29",
          4926 => x"08",
          4927 => x"a0",
          4928 => x"82",
          4929 => x"51",
          4930 => x"d5",
          4931 => x"71",
          4932 => x"c8",
          4933 => x"82",
          4934 => x"a7",
          4935 => x"c8",
          4936 => x"38",
          4937 => x"08",
          4938 => x"d6",
          4939 => x"0b",
          4940 => x"08",
          4941 => x"98",
          4942 => x"c4",
          4943 => x"82",
          4944 => x"80",
          4945 => x"d8",
          4946 => x"0d",
          4947 => x"82",
          4948 => x"04",
          4949 => x"83",
          4950 => x"82",
          4951 => x"84",
          4952 => x"d6",
          4953 => x"80",
          4954 => x"83",
          4955 => x"ff",
          4956 => x"82",
          4957 => x"54",
          4958 => x"74",
          4959 => x"76",
          4960 => x"82",
          4961 => x"54",
          4962 => x"34",
          4963 => x"34",
          4964 => x"08",
          4965 => x"15",
          4966 => x"15",
          4967 => x"d0",
          4968 => x"cc",
          4969 => x"fe",
          4970 => x"70",
          4971 => x"06",
          4972 => x"58",
          4973 => x"74",
          4974 => x"73",
          4975 => x"82",
          4976 => x"70",
          4977 => x"d6",
          4978 => x"f8",
          4979 => x"55",
          4980 => x"34",
          4981 => x"34",
          4982 => x"04",
          4983 => x"73",
          4984 => x"84",
          4985 => x"38",
          4986 => x"2a",
          4987 => x"83",
          4988 => x"51",
          4989 => x"82",
          4990 => x"83",
          4991 => x"f9",
          4992 => x"a6",
          4993 => x"84",
          4994 => x"22",
          4995 => x"d6",
          4996 => x"83",
          4997 => x"74",
          4998 => x"11",
          4999 => x"12",
          5000 => x"2b",
          5001 => x"05",
          5002 => x"71",
          5003 => x"06",
          5004 => x"2a",
          5005 => x"59",
          5006 => x"57",
          5007 => x"71",
          5008 => x"81",
          5009 => x"d6",
          5010 => x"75",
          5011 => x"54",
          5012 => x"34",
          5013 => x"34",
          5014 => x"08",
          5015 => x"33",
          5016 => x"71",
          5017 => x"70",
          5018 => x"ff",
          5019 => x"52",
          5020 => x"05",
          5021 => x"ff",
          5022 => x"2a",
          5023 => x"71",
          5024 => x"72",
          5025 => x"53",
          5026 => x"34",
          5027 => x"08",
          5028 => x"76",
          5029 => x"17",
          5030 => x"0d",
          5031 => x"0d",
          5032 => x"08",
          5033 => x"9e",
          5034 => x"83",
          5035 => x"86",
          5036 => x"12",
          5037 => x"2b",
          5038 => x"07",
          5039 => x"52",
          5040 => x"05",
          5041 => x"85",
          5042 => x"88",
          5043 => x"88",
          5044 => x"56",
          5045 => x"13",
          5046 => x"13",
          5047 => x"d0",
          5048 => x"84",
          5049 => x"12",
          5050 => x"2b",
          5051 => x"07",
          5052 => x"52",
          5053 => x"12",
          5054 => x"33",
          5055 => x"07",
          5056 => x"54",
          5057 => x"70",
          5058 => x"73",
          5059 => x"82",
          5060 => x"13",
          5061 => x"12",
          5062 => x"2b",
          5063 => x"ff",
          5064 => x"88",
          5065 => x"53",
          5066 => x"73",
          5067 => x"14",
          5068 => x"0d",
          5069 => x"0d",
          5070 => x"22",
          5071 => x"08",
          5072 => x"71",
          5073 => x"81",
          5074 => x"88",
          5075 => x"88",
          5076 => x"33",
          5077 => x"71",
          5078 => x"90",
          5079 => x"5f",
          5080 => x"5a",
          5081 => x"54",
          5082 => x"80",
          5083 => x"51",
          5084 => x"82",
          5085 => x"70",
          5086 => x"81",
          5087 => x"8b",
          5088 => x"2b",
          5089 => x"70",
          5090 => x"33",
          5091 => x"07",
          5092 => x"8f",
          5093 => x"51",
          5094 => x"53",
          5095 => x"72",
          5096 => x"2a",
          5097 => x"82",
          5098 => x"83",
          5099 => x"d6",
          5100 => x"16",
          5101 => x"12",
          5102 => x"2b",
          5103 => x"07",
          5104 => x"55",
          5105 => x"33",
          5106 => x"71",
          5107 => x"70",
          5108 => x"06",
          5109 => x"57",
          5110 => x"52",
          5111 => x"71",
          5112 => x"88",
          5113 => x"fb",
          5114 => x"d6",
          5115 => x"84",
          5116 => x"22",
          5117 => x"72",
          5118 => x"33",
          5119 => x"71",
          5120 => x"83",
          5121 => x"5b",
          5122 => x"52",
          5123 => x"33",
          5124 => x"71",
          5125 => x"02",
          5126 => x"05",
          5127 => x"70",
          5128 => x"51",
          5129 => x"71",
          5130 => x"81",
          5131 => x"d6",
          5132 => x"15",
          5133 => x"12",
          5134 => x"2b",
          5135 => x"07",
          5136 => x"52",
          5137 => x"12",
          5138 => x"33",
          5139 => x"07",
          5140 => x"54",
          5141 => x"70",
          5142 => x"72",
          5143 => x"82",
          5144 => x"14",
          5145 => x"83",
          5146 => x"88",
          5147 => x"d6",
          5148 => x"54",
          5149 => x"04",
          5150 => x"7b",
          5151 => x"08",
          5152 => x"70",
          5153 => x"06",
          5154 => x"53",
          5155 => x"82",
          5156 => x"76",
          5157 => x"11",
          5158 => x"83",
          5159 => x"8b",
          5160 => x"2b",
          5161 => x"70",
          5162 => x"33",
          5163 => x"71",
          5164 => x"53",
          5165 => x"53",
          5166 => x"59",
          5167 => x"25",
          5168 => x"80",
          5169 => x"51",
          5170 => x"81",
          5171 => x"14",
          5172 => x"33",
          5173 => x"71",
          5174 => x"76",
          5175 => x"2a",
          5176 => x"58",
          5177 => x"14",
          5178 => x"ff",
          5179 => x"87",
          5180 => x"d6",
          5181 => x"19",
          5182 => x"85",
          5183 => x"88",
          5184 => x"88",
          5185 => x"5b",
          5186 => x"84",
          5187 => x"85",
          5188 => x"d6",
          5189 => x"53",
          5190 => x"14",
          5191 => x"87",
          5192 => x"d6",
          5193 => x"76",
          5194 => x"75",
          5195 => x"82",
          5196 => x"18",
          5197 => x"12",
          5198 => x"2b",
          5199 => x"80",
          5200 => x"88",
          5201 => x"55",
          5202 => x"74",
          5203 => x"15",
          5204 => x"0d",
          5205 => x"0d",
          5206 => x"d6",
          5207 => x"38",
          5208 => x"71",
          5209 => x"38",
          5210 => x"8c",
          5211 => x"0d",
          5212 => x"0d",
          5213 => x"58",
          5214 => x"82",
          5215 => x"83",
          5216 => x"82",
          5217 => x"84",
          5218 => x"12",
          5219 => x"2b",
          5220 => x"59",
          5221 => x"81",
          5222 => x"75",
          5223 => x"cb",
          5224 => x"29",
          5225 => x"81",
          5226 => x"88",
          5227 => x"81",
          5228 => x"79",
          5229 => x"ff",
          5230 => x"7f",
          5231 => x"51",
          5232 => x"77",
          5233 => x"38",
          5234 => x"85",
          5235 => x"5a",
          5236 => x"33",
          5237 => x"71",
          5238 => x"57",
          5239 => x"38",
          5240 => x"ff",
          5241 => x"7a",
          5242 => x"80",
          5243 => x"82",
          5244 => x"11",
          5245 => x"12",
          5246 => x"2b",
          5247 => x"ff",
          5248 => x"52",
          5249 => x"55",
          5250 => x"83",
          5251 => x"80",
          5252 => x"26",
          5253 => x"74",
          5254 => x"2e",
          5255 => x"77",
          5256 => x"81",
          5257 => x"75",
          5258 => x"3f",
          5259 => x"82",
          5260 => x"79",
          5261 => x"f7",
          5262 => x"d6",
          5263 => x"1c",
          5264 => x"87",
          5265 => x"8b",
          5266 => x"2b",
          5267 => x"5e",
          5268 => x"7a",
          5269 => x"ff",
          5270 => x"88",
          5271 => x"56",
          5272 => x"15",
          5273 => x"ff",
          5274 => x"85",
          5275 => x"d6",
          5276 => x"83",
          5277 => x"72",
          5278 => x"33",
          5279 => x"71",
          5280 => x"70",
          5281 => x"5b",
          5282 => x"56",
          5283 => x"19",
          5284 => x"19",
          5285 => x"d0",
          5286 => x"84",
          5287 => x"12",
          5288 => x"2b",
          5289 => x"07",
          5290 => x"55",
          5291 => x"78",
          5292 => x"76",
          5293 => x"82",
          5294 => x"70",
          5295 => x"84",
          5296 => x"12",
          5297 => x"2b",
          5298 => x"2a",
          5299 => x"52",
          5300 => x"84",
          5301 => x"85",
          5302 => x"d6",
          5303 => x"84",
          5304 => x"82",
          5305 => x"8d",
          5306 => x"fe",
          5307 => x"52",
          5308 => x"08",
          5309 => x"dc",
          5310 => x"71",
          5311 => x"38",
          5312 => x"ed",
          5313 => x"d8",
          5314 => x"82",
          5315 => x"84",
          5316 => x"ee",
          5317 => x"66",
          5318 => x"70",
          5319 => x"d6",
          5320 => x"2e",
          5321 => x"84",
          5322 => x"3f",
          5323 => x"7e",
          5324 => x"3f",
          5325 => x"08",
          5326 => x"39",
          5327 => x"7b",
          5328 => x"3f",
          5329 => x"ba",
          5330 => x"f5",
          5331 => x"d6",
          5332 => x"ff",
          5333 => x"d6",
          5334 => x"71",
          5335 => x"70",
          5336 => x"06",
          5337 => x"73",
          5338 => x"81",
          5339 => x"88",
          5340 => x"75",
          5341 => x"ff",
          5342 => x"88",
          5343 => x"73",
          5344 => x"70",
          5345 => x"33",
          5346 => x"07",
          5347 => x"53",
          5348 => x"48",
          5349 => x"54",
          5350 => x"56",
          5351 => x"80",
          5352 => x"76",
          5353 => x"06",
          5354 => x"83",
          5355 => x"42",
          5356 => x"33",
          5357 => x"71",
          5358 => x"70",
          5359 => x"70",
          5360 => x"33",
          5361 => x"71",
          5362 => x"53",
          5363 => x"56",
          5364 => x"25",
          5365 => x"75",
          5366 => x"ff",
          5367 => x"54",
          5368 => x"81",
          5369 => x"18",
          5370 => x"2e",
          5371 => x"8f",
          5372 => x"f6",
          5373 => x"83",
          5374 => x"58",
          5375 => x"7f",
          5376 => x"74",
          5377 => x"78",
          5378 => x"3f",
          5379 => x"7f",
          5380 => x"75",
          5381 => x"38",
          5382 => x"11",
          5383 => x"33",
          5384 => x"07",
          5385 => x"f4",
          5386 => x"52",
          5387 => x"b7",
          5388 => x"d8",
          5389 => x"ff",
          5390 => x"7c",
          5391 => x"2b",
          5392 => x"08",
          5393 => x"53",
          5394 => x"90",
          5395 => x"d6",
          5396 => x"84",
          5397 => x"ff",
          5398 => x"5c",
          5399 => x"60",
          5400 => x"74",
          5401 => x"38",
          5402 => x"c9",
          5403 => x"d0",
          5404 => x"11",
          5405 => x"33",
          5406 => x"07",
          5407 => x"f4",
          5408 => x"52",
          5409 => x"df",
          5410 => x"d8",
          5411 => x"ff",
          5412 => x"7c",
          5413 => x"2b",
          5414 => x"08",
          5415 => x"53",
          5416 => x"8f",
          5417 => x"d6",
          5418 => x"84",
          5419 => x"05",
          5420 => x"73",
          5421 => x"06",
          5422 => x"7b",
          5423 => x"f9",
          5424 => x"d6",
          5425 => x"82",
          5426 => x"80",
          5427 => x"7d",
          5428 => x"82",
          5429 => x"51",
          5430 => x"3f",
          5431 => x"98",
          5432 => x"7a",
          5433 => x"38",
          5434 => x"52",
          5435 => x"8f",
          5436 => x"83",
          5437 => x"d0",
          5438 => x"05",
          5439 => x"3f",
          5440 => x"82",
          5441 => x"94",
          5442 => x"fc",
          5443 => x"77",
          5444 => x"54",
          5445 => x"82",
          5446 => x"55",
          5447 => x"08",
          5448 => x"38",
          5449 => x"52",
          5450 => x"08",
          5451 => x"e4",
          5452 => x"d6",
          5453 => x"3d",
          5454 => x"3d",
          5455 => x"05",
          5456 => x"52",
          5457 => x"87",
          5458 => x"d4",
          5459 => x"71",
          5460 => x"0c",
          5461 => x"04",
          5462 => x"02",
          5463 => x"02",
          5464 => x"05",
          5465 => x"83",
          5466 => x"26",
          5467 => x"72",
          5468 => x"c0",
          5469 => x"53",
          5470 => x"74",
          5471 => x"38",
          5472 => x"73",
          5473 => x"c0",
          5474 => x"51",
          5475 => x"85",
          5476 => x"98",
          5477 => x"52",
          5478 => x"82",
          5479 => x"70",
          5480 => x"38",
          5481 => x"8c",
          5482 => x"ec",
          5483 => x"fc",
          5484 => x"52",
          5485 => x"87",
          5486 => x"08",
          5487 => x"2e",
          5488 => x"82",
          5489 => x"34",
          5490 => x"13",
          5491 => x"82",
          5492 => x"86",
          5493 => x"f3",
          5494 => x"62",
          5495 => x"05",
          5496 => x"57",
          5497 => x"83",
          5498 => x"fe",
          5499 => x"d6",
          5500 => x"06",
          5501 => x"71",
          5502 => x"71",
          5503 => x"2b",
          5504 => x"80",
          5505 => x"92",
          5506 => x"c0",
          5507 => x"41",
          5508 => x"5a",
          5509 => x"87",
          5510 => x"0c",
          5511 => x"84",
          5512 => x"08",
          5513 => x"70",
          5514 => x"53",
          5515 => x"2e",
          5516 => x"08",
          5517 => x"70",
          5518 => x"34",
          5519 => x"80",
          5520 => x"53",
          5521 => x"2e",
          5522 => x"53",
          5523 => x"26",
          5524 => x"80",
          5525 => x"87",
          5526 => x"08",
          5527 => x"38",
          5528 => x"8c",
          5529 => x"80",
          5530 => x"78",
          5531 => x"99",
          5532 => x"0c",
          5533 => x"8c",
          5534 => x"08",
          5535 => x"51",
          5536 => x"38",
          5537 => x"8d",
          5538 => x"17",
          5539 => x"81",
          5540 => x"53",
          5541 => x"2e",
          5542 => x"fc",
          5543 => x"52",
          5544 => x"7d",
          5545 => x"ed",
          5546 => x"80",
          5547 => x"71",
          5548 => x"38",
          5549 => x"53",
          5550 => x"d8",
          5551 => x"0d",
          5552 => x"0d",
          5553 => x"02",
          5554 => x"05",
          5555 => x"58",
          5556 => x"80",
          5557 => x"fc",
          5558 => x"d6",
          5559 => x"06",
          5560 => x"71",
          5561 => x"81",
          5562 => x"38",
          5563 => x"2b",
          5564 => x"80",
          5565 => x"92",
          5566 => x"c0",
          5567 => x"40",
          5568 => x"5a",
          5569 => x"c0",
          5570 => x"76",
          5571 => x"76",
          5572 => x"75",
          5573 => x"2a",
          5574 => x"51",
          5575 => x"80",
          5576 => x"7a",
          5577 => x"5c",
          5578 => x"81",
          5579 => x"81",
          5580 => x"06",
          5581 => x"80",
          5582 => x"87",
          5583 => x"08",
          5584 => x"38",
          5585 => x"8c",
          5586 => x"80",
          5587 => x"77",
          5588 => x"99",
          5589 => x"0c",
          5590 => x"8c",
          5591 => x"08",
          5592 => x"51",
          5593 => x"38",
          5594 => x"8d",
          5595 => x"70",
          5596 => x"84",
          5597 => x"5b",
          5598 => x"2e",
          5599 => x"fc",
          5600 => x"52",
          5601 => x"7d",
          5602 => x"f8",
          5603 => x"80",
          5604 => x"71",
          5605 => x"38",
          5606 => x"53",
          5607 => x"d8",
          5608 => x"0d",
          5609 => x"0d",
          5610 => x"05",
          5611 => x"02",
          5612 => x"05",
          5613 => x"54",
          5614 => x"fe",
          5615 => x"d8",
          5616 => x"53",
          5617 => x"80",
          5618 => x"0b",
          5619 => x"8c",
          5620 => x"71",
          5621 => x"dc",
          5622 => x"24",
          5623 => x"84",
          5624 => x"92",
          5625 => x"54",
          5626 => x"8d",
          5627 => x"39",
          5628 => x"80",
          5629 => x"cb",
          5630 => x"70",
          5631 => x"81",
          5632 => x"52",
          5633 => x"8a",
          5634 => x"98",
          5635 => x"71",
          5636 => x"c0",
          5637 => x"52",
          5638 => x"81",
          5639 => x"c0",
          5640 => x"53",
          5641 => x"82",
          5642 => x"71",
          5643 => x"39",
          5644 => x"39",
          5645 => x"77",
          5646 => x"81",
          5647 => x"72",
          5648 => x"84",
          5649 => x"73",
          5650 => x"0c",
          5651 => x"04",
          5652 => x"74",
          5653 => x"71",
          5654 => x"2b",
          5655 => x"d8",
          5656 => x"84",
          5657 => x"fd",
          5658 => x"83",
          5659 => x"12",
          5660 => x"2b",
          5661 => x"07",
          5662 => x"70",
          5663 => x"2b",
          5664 => x"07",
          5665 => x"0c",
          5666 => x"56",
          5667 => x"3d",
          5668 => x"3d",
          5669 => x"84",
          5670 => x"22",
          5671 => x"72",
          5672 => x"54",
          5673 => x"2a",
          5674 => x"34",
          5675 => x"04",
          5676 => x"73",
          5677 => x"70",
          5678 => x"05",
          5679 => x"88",
          5680 => x"72",
          5681 => x"54",
          5682 => x"2a",
          5683 => x"70",
          5684 => x"34",
          5685 => x"51",
          5686 => x"83",
          5687 => x"fe",
          5688 => x"75",
          5689 => x"51",
          5690 => x"92",
          5691 => x"81",
          5692 => x"73",
          5693 => x"55",
          5694 => x"51",
          5695 => x"3d",
          5696 => x"3d",
          5697 => x"76",
          5698 => x"72",
          5699 => x"05",
          5700 => x"11",
          5701 => x"38",
          5702 => x"04",
          5703 => x"78",
          5704 => x"56",
          5705 => x"81",
          5706 => x"74",
          5707 => x"56",
          5708 => x"31",
          5709 => x"52",
          5710 => x"80",
          5711 => x"71",
          5712 => x"38",
          5713 => x"d8",
          5714 => x"0d",
          5715 => x"0d",
          5716 => x"51",
          5717 => x"73",
          5718 => x"81",
          5719 => x"33",
          5720 => x"38",
          5721 => x"d6",
          5722 => x"3d",
          5723 => x"0b",
          5724 => x"0c",
          5725 => x"0d",
          5726 => x"70",
          5727 => x"52",
          5728 => x"55",
          5729 => x"3f",
          5730 => x"d6",
          5731 => x"38",
          5732 => x"98",
          5733 => x"52",
          5734 => x"f7",
          5735 => x"d6",
          5736 => x"ff",
          5737 => x"72",
          5738 => x"38",
          5739 => x"72",
          5740 => x"d6",
          5741 => x"3d",
          5742 => x"3d",
          5743 => x"80",
          5744 => x"33",
          5745 => x"7a",
          5746 => x"38",
          5747 => x"16",
          5748 => x"16",
          5749 => x"17",
          5750 => x"f9",
          5751 => x"d6",
          5752 => x"2e",
          5753 => x"b7",
          5754 => x"d8",
          5755 => x"34",
          5756 => x"70",
          5757 => x"31",
          5758 => x"59",
          5759 => x"77",
          5760 => x"82",
          5761 => x"74",
          5762 => x"81",
          5763 => x"81",
          5764 => x"53",
          5765 => x"16",
          5766 => x"a5",
          5767 => x"81",
          5768 => x"d6",
          5769 => x"3d",
          5770 => x"3d",
          5771 => x"56",
          5772 => x"74",
          5773 => x"2e",
          5774 => x"51",
          5775 => x"82",
          5776 => x"57",
          5777 => x"08",
          5778 => x"54",
          5779 => x"16",
          5780 => x"33",
          5781 => x"3f",
          5782 => x"08",
          5783 => x"38",
          5784 => x"57",
          5785 => x"0c",
          5786 => x"d8",
          5787 => x"0d",
          5788 => x"0d",
          5789 => x"57",
          5790 => x"82",
          5791 => x"58",
          5792 => x"08",
          5793 => x"76",
          5794 => x"83",
          5795 => x"06",
          5796 => x"84",
          5797 => x"78",
          5798 => x"81",
          5799 => x"38",
          5800 => x"82",
          5801 => x"52",
          5802 => x"52",
          5803 => x"3f",
          5804 => x"52",
          5805 => x"51",
          5806 => x"84",
          5807 => x"d2",
          5808 => x"fb",
          5809 => x"8a",
          5810 => x"52",
          5811 => x"51",
          5812 => x"94",
          5813 => x"84",
          5814 => x"fb",
          5815 => x"17",
          5816 => x"a4",
          5817 => x"c8",
          5818 => x"08",
          5819 => x"b4",
          5820 => x"55",
          5821 => x"81",
          5822 => x"f7",
          5823 => x"84",
          5824 => x"53",
          5825 => x"17",
          5826 => x"99",
          5827 => x"d8",
          5828 => x"83",
          5829 => x"77",
          5830 => x"0c",
          5831 => x"04",
          5832 => x"77",
          5833 => x"12",
          5834 => x"55",
          5835 => x"56",
          5836 => x"8d",
          5837 => x"22",
          5838 => x"b0",
          5839 => x"57",
          5840 => x"d6",
          5841 => x"3d",
          5842 => x"3d",
          5843 => x"70",
          5844 => x"57",
          5845 => x"81",
          5846 => x"9c",
          5847 => x"81",
          5848 => x"74",
          5849 => x"72",
          5850 => x"f5",
          5851 => x"24",
          5852 => x"81",
          5853 => x"81",
          5854 => x"83",
          5855 => x"38",
          5856 => x"76",
          5857 => x"70",
          5858 => x"16",
          5859 => x"74",
          5860 => x"96",
          5861 => x"d8",
          5862 => x"38",
          5863 => x"06",
          5864 => x"33",
          5865 => x"89",
          5866 => x"08",
          5867 => x"54",
          5868 => x"fc",
          5869 => x"d6",
          5870 => x"fe",
          5871 => x"ff",
          5872 => x"11",
          5873 => x"2b",
          5874 => x"81",
          5875 => x"2a",
          5876 => x"51",
          5877 => x"e2",
          5878 => x"ff",
          5879 => x"da",
          5880 => x"2a",
          5881 => x"05",
          5882 => x"fc",
          5883 => x"d6",
          5884 => x"c6",
          5885 => x"83",
          5886 => x"05",
          5887 => x"f8",
          5888 => x"d6",
          5889 => x"ff",
          5890 => x"ae",
          5891 => x"2a",
          5892 => x"05",
          5893 => x"fc",
          5894 => x"d6",
          5895 => x"38",
          5896 => x"83",
          5897 => x"05",
          5898 => x"f8",
          5899 => x"d6",
          5900 => x"0a",
          5901 => x"39",
          5902 => x"82",
          5903 => x"89",
          5904 => x"f8",
          5905 => x"7c",
          5906 => x"56",
          5907 => x"77",
          5908 => x"38",
          5909 => x"08",
          5910 => x"38",
          5911 => x"72",
          5912 => x"9d",
          5913 => x"24",
          5914 => x"81",
          5915 => x"82",
          5916 => x"83",
          5917 => x"38",
          5918 => x"76",
          5919 => x"70",
          5920 => x"18",
          5921 => x"76",
          5922 => x"9e",
          5923 => x"d8",
          5924 => x"d6",
          5925 => x"d9",
          5926 => x"ff",
          5927 => x"05",
          5928 => x"81",
          5929 => x"54",
          5930 => x"80",
          5931 => x"77",
          5932 => x"f0",
          5933 => x"8f",
          5934 => x"51",
          5935 => x"34",
          5936 => x"17",
          5937 => x"2a",
          5938 => x"05",
          5939 => x"fa",
          5940 => x"d6",
          5941 => x"82",
          5942 => x"81",
          5943 => x"83",
          5944 => x"b8",
          5945 => x"2a",
          5946 => x"8f",
          5947 => x"2a",
          5948 => x"f0",
          5949 => x"06",
          5950 => x"72",
          5951 => x"ec",
          5952 => x"2a",
          5953 => x"05",
          5954 => x"fa",
          5955 => x"d6",
          5956 => x"82",
          5957 => x"80",
          5958 => x"83",
          5959 => x"52",
          5960 => x"fe",
          5961 => x"b8",
          5962 => x"e6",
          5963 => x"76",
          5964 => x"17",
          5965 => x"75",
          5966 => x"3f",
          5967 => x"08",
          5968 => x"d8",
          5969 => x"77",
          5970 => x"77",
          5971 => x"fc",
          5972 => x"b8",
          5973 => x"51",
          5974 => x"8b",
          5975 => x"d8",
          5976 => x"06",
          5977 => x"72",
          5978 => x"3f",
          5979 => x"17",
          5980 => x"d6",
          5981 => x"3d",
          5982 => x"3d",
          5983 => x"7e",
          5984 => x"56",
          5985 => x"75",
          5986 => x"74",
          5987 => x"27",
          5988 => x"80",
          5989 => x"ff",
          5990 => x"75",
          5991 => x"3f",
          5992 => x"08",
          5993 => x"d8",
          5994 => x"38",
          5995 => x"54",
          5996 => x"81",
          5997 => x"39",
          5998 => x"08",
          5999 => x"39",
          6000 => x"51",
          6001 => x"82",
          6002 => x"58",
          6003 => x"08",
          6004 => x"c7",
          6005 => x"d8",
          6006 => x"d2",
          6007 => x"d8",
          6008 => x"cf",
          6009 => x"74",
          6010 => x"fc",
          6011 => x"d6",
          6012 => x"38",
          6013 => x"fe",
          6014 => x"08",
          6015 => x"74",
          6016 => x"38",
          6017 => x"17",
          6018 => x"33",
          6019 => x"73",
          6020 => x"77",
          6021 => x"26",
          6022 => x"80",
          6023 => x"d6",
          6024 => x"3d",
          6025 => x"3d",
          6026 => x"71",
          6027 => x"5b",
          6028 => x"90",
          6029 => x"77",
          6030 => x"38",
          6031 => x"78",
          6032 => x"81",
          6033 => x"79",
          6034 => x"f9",
          6035 => x"55",
          6036 => x"d8",
          6037 => x"e0",
          6038 => x"d8",
          6039 => x"d6",
          6040 => x"2e",
          6041 => x"9c",
          6042 => x"d6",
          6043 => x"82",
          6044 => x"58",
          6045 => x"70",
          6046 => x"80",
          6047 => x"38",
          6048 => x"09",
          6049 => x"e2",
          6050 => x"56",
          6051 => x"76",
          6052 => x"82",
          6053 => x"7a",
          6054 => x"3f",
          6055 => x"d6",
          6056 => x"2e",
          6057 => x"86",
          6058 => x"d8",
          6059 => x"d6",
          6060 => x"70",
          6061 => x"07",
          6062 => x"7c",
          6063 => x"d8",
          6064 => x"51",
          6065 => x"81",
          6066 => x"d6",
          6067 => x"2e",
          6068 => x"17",
          6069 => x"74",
          6070 => x"73",
          6071 => x"27",
          6072 => x"58",
          6073 => x"80",
          6074 => x"56",
          6075 => x"9c",
          6076 => x"26",
          6077 => x"56",
          6078 => x"81",
          6079 => x"52",
          6080 => x"c6",
          6081 => x"d8",
          6082 => x"b8",
          6083 => x"82",
          6084 => x"81",
          6085 => x"06",
          6086 => x"d6",
          6087 => x"82",
          6088 => x"09",
          6089 => x"72",
          6090 => x"70",
          6091 => x"51",
          6092 => x"80",
          6093 => x"78",
          6094 => x"06",
          6095 => x"73",
          6096 => x"39",
          6097 => x"52",
          6098 => x"f7",
          6099 => x"d8",
          6100 => x"d8",
          6101 => x"82",
          6102 => x"07",
          6103 => x"55",
          6104 => x"2e",
          6105 => x"80",
          6106 => x"75",
          6107 => x"76",
          6108 => x"3f",
          6109 => x"08",
          6110 => x"38",
          6111 => x"0c",
          6112 => x"fe",
          6113 => x"08",
          6114 => x"74",
          6115 => x"ff",
          6116 => x"0c",
          6117 => x"81",
          6118 => x"84",
          6119 => x"39",
          6120 => x"81",
          6121 => x"8c",
          6122 => x"8c",
          6123 => x"d8",
          6124 => x"39",
          6125 => x"55",
          6126 => x"d8",
          6127 => x"0d",
          6128 => x"0d",
          6129 => x"55",
          6130 => x"82",
          6131 => x"58",
          6132 => x"d6",
          6133 => x"d8",
          6134 => x"74",
          6135 => x"3f",
          6136 => x"08",
          6137 => x"08",
          6138 => x"59",
          6139 => x"77",
          6140 => x"70",
          6141 => x"8a",
          6142 => x"84",
          6143 => x"56",
          6144 => x"58",
          6145 => x"97",
          6146 => x"75",
          6147 => x"52",
          6148 => x"51",
          6149 => x"82",
          6150 => x"80",
          6151 => x"8a",
          6152 => x"32",
          6153 => x"72",
          6154 => x"2a",
          6155 => x"56",
          6156 => x"d8",
          6157 => x"0d",
          6158 => x"0d",
          6159 => x"08",
          6160 => x"74",
          6161 => x"26",
          6162 => x"74",
          6163 => x"72",
          6164 => x"74",
          6165 => x"88",
          6166 => x"73",
          6167 => x"33",
          6168 => x"27",
          6169 => x"16",
          6170 => x"9b",
          6171 => x"2a",
          6172 => x"88",
          6173 => x"58",
          6174 => x"80",
          6175 => x"16",
          6176 => x"0c",
          6177 => x"8a",
          6178 => x"89",
          6179 => x"72",
          6180 => x"38",
          6181 => x"51",
          6182 => x"82",
          6183 => x"54",
          6184 => x"08",
          6185 => x"38",
          6186 => x"d6",
          6187 => x"8b",
          6188 => x"08",
          6189 => x"08",
          6190 => x"82",
          6191 => x"74",
          6192 => x"cb",
          6193 => x"75",
          6194 => x"3f",
          6195 => x"08",
          6196 => x"73",
          6197 => x"98",
          6198 => x"82",
          6199 => x"2e",
          6200 => x"39",
          6201 => x"39",
          6202 => x"13",
          6203 => x"74",
          6204 => x"16",
          6205 => x"18",
          6206 => x"77",
          6207 => x"0c",
          6208 => x"04",
          6209 => x"7a",
          6210 => x"12",
          6211 => x"59",
          6212 => x"80",
          6213 => x"86",
          6214 => x"98",
          6215 => x"14",
          6216 => x"55",
          6217 => x"81",
          6218 => x"83",
          6219 => x"77",
          6220 => x"81",
          6221 => x"0c",
          6222 => x"55",
          6223 => x"76",
          6224 => x"17",
          6225 => x"74",
          6226 => x"9b",
          6227 => x"39",
          6228 => x"ff",
          6229 => x"2a",
          6230 => x"81",
          6231 => x"52",
          6232 => x"e6",
          6233 => x"d8",
          6234 => x"55",
          6235 => x"d6",
          6236 => x"80",
          6237 => x"55",
          6238 => x"08",
          6239 => x"f4",
          6240 => x"08",
          6241 => x"08",
          6242 => x"38",
          6243 => x"77",
          6244 => x"84",
          6245 => x"39",
          6246 => x"52",
          6247 => x"86",
          6248 => x"d8",
          6249 => x"55",
          6250 => x"08",
          6251 => x"c4",
          6252 => x"82",
          6253 => x"81",
          6254 => x"81",
          6255 => x"d8",
          6256 => x"b0",
          6257 => x"d8",
          6258 => x"51",
          6259 => x"82",
          6260 => x"a0",
          6261 => x"15",
          6262 => x"75",
          6263 => x"3f",
          6264 => x"08",
          6265 => x"76",
          6266 => x"77",
          6267 => x"9c",
          6268 => x"55",
          6269 => x"d8",
          6270 => x"0d",
          6271 => x"0d",
          6272 => x"08",
          6273 => x"80",
          6274 => x"fc",
          6275 => x"d6",
          6276 => x"82",
          6277 => x"80",
          6278 => x"d6",
          6279 => x"98",
          6280 => x"78",
          6281 => x"3f",
          6282 => x"08",
          6283 => x"d8",
          6284 => x"38",
          6285 => x"08",
          6286 => x"70",
          6287 => x"58",
          6288 => x"2e",
          6289 => x"83",
          6290 => x"82",
          6291 => x"55",
          6292 => x"81",
          6293 => x"07",
          6294 => x"2e",
          6295 => x"16",
          6296 => x"2e",
          6297 => x"88",
          6298 => x"82",
          6299 => x"56",
          6300 => x"51",
          6301 => x"82",
          6302 => x"54",
          6303 => x"08",
          6304 => x"9b",
          6305 => x"2e",
          6306 => x"83",
          6307 => x"73",
          6308 => x"0c",
          6309 => x"04",
          6310 => x"76",
          6311 => x"54",
          6312 => x"82",
          6313 => x"83",
          6314 => x"76",
          6315 => x"53",
          6316 => x"2e",
          6317 => x"90",
          6318 => x"51",
          6319 => x"82",
          6320 => x"90",
          6321 => x"53",
          6322 => x"d8",
          6323 => x"0d",
          6324 => x"0d",
          6325 => x"83",
          6326 => x"54",
          6327 => x"55",
          6328 => x"3f",
          6329 => x"51",
          6330 => x"2e",
          6331 => x"8b",
          6332 => x"2a",
          6333 => x"51",
          6334 => x"86",
          6335 => x"fd",
          6336 => x"54",
          6337 => x"53",
          6338 => x"71",
          6339 => x"05",
          6340 => x"05",
          6341 => x"05",
          6342 => x"06",
          6343 => x"51",
          6344 => x"e4",
          6345 => x"d6",
          6346 => x"3d",
          6347 => x"3d",
          6348 => x"40",
          6349 => x"08",
          6350 => x"ff",
          6351 => x"98",
          6352 => x"2e",
          6353 => x"98",
          6354 => x"7d",
          6355 => x"3f",
          6356 => x"08",
          6357 => x"d8",
          6358 => x"38",
          6359 => x"70",
          6360 => x"73",
          6361 => x"5b",
          6362 => x"8b",
          6363 => x"06",
          6364 => x"06",
          6365 => x"86",
          6366 => x"d6",
          6367 => x"73",
          6368 => x"09",
          6369 => x"38",
          6370 => x"d6",
          6371 => x"73",
          6372 => x"81",
          6373 => x"81",
          6374 => x"07",
          6375 => x"38",
          6376 => x"08",
          6377 => x"54",
          6378 => x"2e",
          6379 => x"83",
          6380 => x"75",
          6381 => x"38",
          6382 => x"81",
          6383 => x"8f",
          6384 => x"06",
          6385 => x"73",
          6386 => x"81",
          6387 => x"72",
          6388 => x"38",
          6389 => x"74",
          6390 => x"70",
          6391 => x"ac",
          6392 => x"5d",
          6393 => x"2e",
          6394 => x"81",
          6395 => x"15",
          6396 => x"73",
          6397 => x"06",
          6398 => x"8c",
          6399 => x"16",
          6400 => x"cc",
          6401 => x"d8",
          6402 => x"ff",
          6403 => x"80",
          6404 => x"33",
          6405 => x"06",
          6406 => x"05",
          6407 => x"7b",
          6408 => x"c7",
          6409 => x"75",
          6410 => x"a4",
          6411 => x"d8",
          6412 => x"ff",
          6413 => x"80",
          6414 => x"73",
          6415 => x"80",
          6416 => x"10",
          6417 => x"53",
          6418 => x"81",
          6419 => x"39",
          6420 => x"ff",
          6421 => x"06",
          6422 => x"17",
          6423 => x"27",
          6424 => x"33",
          6425 => x"70",
          6426 => x"54",
          6427 => x"2e",
          6428 => x"81",
          6429 => x"38",
          6430 => x"53",
          6431 => x"ff",
          6432 => x"ff",
          6433 => x"84",
          6434 => x"53",
          6435 => x"39",
          6436 => x"74",
          6437 => x"3f",
          6438 => x"08",
          6439 => x"53",
          6440 => x"a7",
          6441 => x"ac",
          6442 => x"39",
          6443 => x"51",
          6444 => x"82",
          6445 => x"5b",
          6446 => x"08",
          6447 => x"19",
          6448 => x"38",
          6449 => x"0b",
          6450 => x"7a",
          6451 => x"0c",
          6452 => x"04",
          6453 => x"60",
          6454 => x"59",
          6455 => x"51",
          6456 => x"82",
          6457 => x"58",
          6458 => x"08",
          6459 => x"81",
          6460 => x"5c",
          6461 => x"1a",
          6462 => x"08",
          6463 => x"ea",
          6464 => x"d6",
          6465 => x"82",
          6466 => x"83",
          6467 => x"19",
          6468 => x"57",
          6469 => x"38",
          6470 => x"f6",
          6471 => x"33",
          6472 => x"81",
          6473 => x"54",
          6474 => x"34",
          6475 => x"2e",
          6476 => x"74",
          6477 => x"81",
          6478 => x"74",
          6479 => x"38",
          6480 => x"38",
          6481 => x"09",
          6482 => x"f7",
          6483 => x"33",
          6484 => x"70",
          6485 => x"55",
          6486 => x"a1",
          6487 => x"2a",
          6488 => x"51",
          6489 => x"2e",
          6490 => x"17",
          6491 => x"bf",
          6492 => x"1c",
          6493 => x"0c",
          6494 => x"75",
          6495 => x"81",
          6496 => x"38",
          6497 => x"56",
          6498 => x"09",
          6499 => x"ac",
          6500 => x"08",
          6501 => x"5d",
          6502 => x"82",
          6503 => x"83",
          6504 => x"55",
          6505 => x"38",
          6506 => x"bf",
          6507 => x"f3",
          6508 => x"81",
          6509 => x"82",
          6510 => x"33",
          6511 => x"e5",
          6512 => x"d6",
          6513 => x"ff",
          6514 => x"79",
          6515 => x"38",
          6516 => x"26",
          6517 => x"75",
          6518 => x"b4",
          6519 => x"d8",
          6520 => x"1e",
          6521 => x"55",
          6522 => x"55",
          6523 => x"3f",
          6524 => x"d8",
          6525 => x"81",
          6526 => x"38",
          6527 => x"39",
          6528 => x"ff",
          6529 => x"06",
          6530 => x"1b",
          6531 => x"27",
          6532 => x"76",
          6533 => x"2a",
          6534 => x"51",
          6535 => x"80",
          6536 => x"73",
          6537 => x"38",
          6538 => x"70",
          6539 => x"73",
          6540 => x"1c",
          6541 => x"06",
          6542 => x"39",
          6543 => x"73",
          6544 => x"7b",
          6545 => x"51",
          6546 => x"82",
          6547 => x"81",
          6548 => x"73",
          6549 => x"38",
          6550 => x"81",
          6551 => x"95",
          6552 => x"a0",
          6553 => x"19",
          6554 => x"b0",
          6555 => x"d8",
          6556 => x"9e",
          6557 => x"5c",
          6558 => x"1a",
          6559 => x"78",
          6560 => x"3f",
          6561 => x"08",
          6562 => x"d8",
          6563 => x"fc",
          6564 => x"82",
          6565 => x"90",
          6566 => x"ee",
          6567 => x"70",
          6568 => x"33",
          6569 => x"56",
          6570 => x"55",
          6571 => x"38",
          6572 => x"08",
          6573 => x"56",
          6574 => x"2e",
          6575 => x"1d",
          6576 => x"70",
          6577 => x"5d",
          6578 => x"53",
          6579 => x"53",
          6580 => x"53",
          6581 => x"87",
          6582 => x"cb",
          6583 => x"06",
          6584 => x"2e",
          6585 => x"80",
          6586 => x"1b",
          6587 => x"8c",
          6588 => x"56",
          6589 => x"7d",
          6590 => x"e3",
          6591 => x"7b",
          6592 => x"38",
          6593 => x"22",
          6594 => x"ff",
          6595 => x"73",
          6596 => x"38",
          6597 => x"ff",
          6598 => x"59",
          6599 => x"74",
          6600 => x"10",
          6601 => x"2a",
          6602 => x"70",
          6603 => x"56",
          6604 => x"80",
          6605 => x"75",
          6606 => x"32",
          6607 => x"57",
          6608 => x"db",
          6609 => x"75",
          6610 => x"84",
          6611 => x"57",
          6612 => x"07",
          6613 => x"b9",
          6614 => x"38",
          6615 => x"73",
          6616 => x"16",
          6617 => x"84",
          6618 => x"56",
          6619 => x"94",
          6620 => x"17",
          6621 => x"74",
          6622 => x"27",
          6623 => x"33",
          6624 => x"2e",
          6625 => x"19",
          6626 => x"54",
          6627 => x"82",
          6628 => x"80",
          6629 => x"ff",
          6630 => x"74",
          6631 => x"81",
          6632 => x"15",
          6633 => x"27",
          6634 => x"19",
          6635 => x"54",
          6636 => x"3d",
          6637 => x"05",
          6638 => x"81",
          6639 => x"a0",
          6640 => x"26",
          6641 => x"17",
          6642 => x"33",
          6643 => x"75",
          6644 => x"75",
          6645 => x"79",
          6646 => x"3f",
          6647 => x"08",
          6648 => x"1b",
          6649 => x"7b",
          6650 => x"38",
          6651 => x"80",
          6652 => x"f0",
          6653 => x"d8",
          6654 => x"d6",
          6655 => x"2e",
          6656 => x"82",
          6657 => x"80",
          6658 => x"ab",
          6659 => x"80",
          6660 => x"70",
          6661 => x"81",
          6662 => x"5e",
          6663 => x"80",
          6664 => x"8d",
          6665 => x"51",
          6666 => x"3f",
          6667 => x"08",
          6668 => x"52",
          6669 => x"c5",
          6670 => x"d8",
          6671 => x"d6",
          6672 => x"9e",
          6673 => x"59",
          6674 => x"81",
          6675 => x"85",
          6676 => x"08",
          6677 => x"54",
          6678 => x"dd",
          6679 => x"d8",
          6680 => x"d6",
          6681 => x"fa",
          6682 => x"51",
          6683 => x"82",
          6684 => x"81",
          6685 => x"98",
          6686 => x"7b",
          6687 => x"3f",
          6688 => x"08",
          6689 => x"d8",
          6690 => x"38",
          6691 => x"9c",
          6692 => x"81",
          6693 => x"57",
          6694 => x"17",
          6695 => x"8b",
          6696 => x"d6",
          6697 => x"17",
          6698 => x"d8",
          6699 => x"16",
          6700 => x"3f",
          6701 => x"f3",
          6702 => x"55",
          6703 => x"ff",
          6704 => x"74",
          6705 => x"22",
          6706 => x"51",
          6707 => x"82",
          6708 => x"33",
          6709 => x"df",
          6710 => x"85",
          6711 => x"ff",
          6712 => x"57",
          6713 => x"d4",
          6714 => x"ff",
          6715 => x"38",
          6716 => x"70",
          6717 => x"73",
          6718 => x"80",
          6719 => x"77",
          6720 => x"0b",
          6721 => x"80",
          6722 => x"ef",
          6723 => x"d6",
          6724 => x"82",
          6725 => x"80",
          6726 => x"19",
          6727 => x"d7",
          6728 => x"08",
          6729 => x"e2",
          6730 => x"d6",
          6731 => x"82",
          6732 => x"ae",
          6733 => x"82",
          6734 => x"52",
          6735 => x"51",
          6736 => x"8b",
          6737 => x"52",
          6738 => x"51",
          6739 => x"9c",
          6740 => x"1b",
          6741 => x"55",
          6742 => x"16",
          6743 => x"83",
          6744 => x"55",
          6745 => x"d8",
          6746 => x"0d",
          6747 => x"0d",
          6748 => x"90",
          6749 => x"13",
          6750 => x"57",
          6751 => x"2e",
          6752 => x"52",
          6753 => x"b1",
          6754 => x"d8",
          6755 => x"d6",
          6756 => x"c9",
          6757 => x"08",
          6758 => x"e1",
          6759 => x"d6",
          6760 => x"82",
          6761 => x"ab",
          6762 => x"08",
          6763 => x"34",
          6764 => x"17",
          6765 => x"08",
          6766 => x"38",
          6767 => x"08",
          6768 => x"ee",
          6769 => x"d6",
          6770 => x"82",
          6771 => x"80",
          6772 => x"73",
          6773 => x"81",
          6774 => x"82",
          6775 => x"d6",
          6776 => x"3d",
          6777 => x"3d",
          6778 => x"71",
          6779 => x"5c",
          6780 => x"19",
          6781 => x"08",
          6782 => x"e2",
          6783 => x"08",
          6784 => x"bb",
          6785 => x"71",
          6786 => x"08",
          6787 => x"57",
          6788 => x"72",
          6789 => x"9d",
          6790 => x"14",
          6791 => x"1b",
          6792 => x"7a",
          6793 => x"d0",
          6794 => x"83",
          6795 => x"51",
          6796 => x"ff",
          6797 => x"74",
          6798 => x"39",
          6799 => x"11",
          6800 => x"31",
          6801 => x"83",
          6802 => x"90",
          6803 => x"51",
          6804 => x"3f",
          6805 => x"08",
          6806 => x"06",
          6807 => x"75",
          6808 => x"81",
          6809 => x"38",
          6810 => x"53",
          6811 => x"74",
          6812 => x"82",
          6813 => x"74",
          6814 => x"70",
          6815 => x"25",
          6816 => x"07",
          6817 => x"73",
          6818 => x"38",
          6819 => x"39",
          6820 => x"81",
          6821 => x"57",
          6822 => x"1d",
          6823 => x"11",
          6824 => x"54",
          6825 => x"f1",
          6826 => x"70",
          6827 => x"30",
          6828 => x"51",
          6829 => x"94",
          6830 => x"0b",
          6831 => x"80",
          6832 => x"58",
          6833 => x"1c",
          6834 => x"33",
          6835 => x"56",
          6836 => x"2e",
          6837 => x"85",
          6838 => x"06",
          6839 => x"e5",
          6840 => x"32",
          6841 => x"72",
          6842 => x"51",
          6843 => x"8b",
          6844 => x"72",
          6845 => x"38",
          6846 => x"81",
          6847 => x"81",
          6848 => x"76",
          6849 => x"58",
          6850 => x"57",
          6851 => x"ff",
          6852 => x"17",
          6853 => x"80",
          6854 => x"34",
          6855 => x"53",
          6856 => x"38",
          6857 => x"bf",
          6858 => x"34",
          6859 => x"e1",
          6860 => x"89",
          6861 => x"5a",
          6862 => x"2e",
          6863 => x"96",
          6864 => x"55",
          6865 => x"ff",
          6866 => x"55",
          6867 => x"aa",
          6868 => x"08",
          6869 => x"51",
          6870 => x"27",
          6871 => x"84",
          6872 => x"39",
          6873 => x"53",
          6874 => x"53",
          6875 => x"8a",
          6876 => x"70",
          6877 => x"06",
          6878 => x"76",
          6879 => x"58",
          6880 => x"81",
          6881 => x"71",
          6882 => x"55",
          6883 => x"b5",
          6884 => x"94",
          6885 => x"0b",
          6886 => x"9c",
          6887 => x"11",
          6888 => x"72",
          6889 => x"89",
          6890 => x"1c",
          6891 => x"13",
          6892 => x"34",
          6893 => x"9c",
          6894 => x"d9",
          6895 => x"d6",
          6896 => x"0c",
          6897 => x"d9",
          6898 => x"d6",
          6899 => x"19",
          6900 => x"51",
          6901 => x"82",
          6902 => x"84",
          6903 => x"3d",
          6904 => x"3d",
          6905 => x"08",
          6906 => x"64",
          6907 => x"55",
          6908 => x"2e",
          6909 => x"55",
          6910 => x"2e",
          6911 => x"80",
          6912 => x"7f",
          6913 => x"88",
          6914 => x"39",
          6915 => x"80",
          6916 => x"56",
          6917 => x"af",
          6918 => x"06",
          6919 => x"56",
          6920 => x"32",
          6921 => x"80",
          6922 => x"51",
          6923 => x"dc",
          6924 => x"1f",
          6925 => x"33",
          6926 => x"9f",
          6927 => x"ff",
          6928 => x"1f",
          6929 => x"7d",
          6930 => x"3f",
          6931 => x"08",
          6932 => x"39",
          6933 => x"08",
          6934 => x"5b",
          6935 => x"92",
          6936 => x"51",
          6937 => x"82",
          6938 => x"ff",
          6939 => x"38",
          6940 => x"0b",
          6941 => x"08",
          6942 => x"78",
          6943 => x"d6",
          6944 => x"2a",
          6945 => x"75",
          6946 => x"59",
          6947 => x"08",
          6948 => x"06",
          6949 => x"70",
          6950 => x"27",
          6951 => x"07",
          6952 => x"56",
          6953 => x"75",
          6954 => x"ae",
          6955 => x"ff",
          6956 => x"75",
          6957 => x"f0",
          6958 => x"3f",
          6959 => x"08",
          6960 => x"78",
          6961 => x"81",
          6962 => x"10",
          6963 => x"74",
          6964 => x"59",
          6965 => x"81",
          6966 => x"61",
          6967 => x"56",
          6968 => x"2e",
          6969 => x"83",
          6970 => x"73",
          6971 => x"70",
          6972 => x"25",
          6973 => x"51",
          6974 => x"38",
          6975 => x"76",
          6976 => x"57",
          6977 => x"09",
          6978 => x"38",
          6979 => x"73",
          6980 => x"38",
          6981 => x"78",
          6982 => x"81",
          6983 => x"38",
          6984 => x"54",
          6985 => x"09",
          6986 => x"c1",
          6987 => x"54",
          6988 => x"09",
          6989 => x"38",
          6990 => x"54",
          6991 => x"80",
          6992 => x"56",
          6993 => x"78",
          6994 => x"38",
          6995 => x"75",
          6996 => x"57",
          6997 => x"58",
          6998 => x"e9",
          6999 => x"07",
          7000 => x"1f",
          7001 => x"39",
          7002 => x"a8",
          7003 => x"1a",
          7004 => x"74",
          7005 => x"71",
          7006 => x"70",
          7007 => x"2a",
          7008 => x"58",
          7009 => x"ae",
          7010 => x"73",
          7011 => x"19",
          7012 => x"38",
          7013 => x"11",
          7014 => x"74",
          7015 => x"38",
          7016 => x"90",
          7017 => x"07",
          7018 => x"39",
          7019 => x"70",
          7020 => x"06",
          7021 => x"73",
          7022 => x"81",
          7023 => x"81",
          7024 => x"1b",
          7025 => x"55",
          7026 => x"2e",
          7027 => x"8f",
          7028 => x"ff",
          7029 => x"73",
          7030 => x"81",
          7031 => x"76",
          7032 => x"78",
          7033 => x"38",
          7034 => x"05",
          7035 => x"54",
          7036 => x"9d",
          7037 => x"1a",
          7038 => x"ff",
          7039 => x"80",
          7040 => x"fe",
          7041 => x"55",
          7042 => x"2e",
          7043 => x"eb",
          7044 => x"a0",
          7045 => x"51",
          7046 => x"80",
          7047 => x"88",
          7048 => x"1a",
          7049 => x"1f",
          7050 => x"75",
          7051 => x"94",
          7052 => x"2e",
          7053 => x"ae",
          7054 => x"70",
          7055 => x"51",
          7056 => x"2e",
          7057 => x"80",
          7058 => x"76",
          7059 => x"d1",
          7060 => x"73",
          7061 => x"26",
          7062 => x"5b",
          7063 => x"70",
          7064 => x"07",
          7065 => x"7e",
          7066 => x"55",
          7067 => x"2e",
          7068 => x"8b",
          7069 => x"38",
          7070 => x"8b",
          7071 => x"07",
          7072 => x"26",
          7073 => x"78",
          7074 => x"8b",
          7075 => x"81",
          7076 => x"5f",
          7077 => x"80",
          7078 => x"af",
          7079 => x"07",
          7080 => x"52",
          7081 => x"cc",
          7082 => x"d6",
          7083 => x"ff",
          7084 => x"87",
          7085 => x"06",
          7086 => x"73",
          7087 => x"38",
          7088 => x"06",
          7089 => x"11",
          7090 => x"81",
          7091 => x"a4",
          7092 => x"54",
          7093 => x"8a",
          7094 => x"07",
          7095 => x"fe",
          7096 => x"18",
          7097 => x"88",
          7098 => x"73",
          7099 => x"18",
          7100 => x"39",
          7101 => x"92",
          7102 => x"82",
          7103 => x"d4",
          7104 => x"d6",
          7105 => x"2e",
          7106 => x"df",
          7107 => x"58",
          7108 => x"ff",
          7109 => x"73",
          7110 => x"38",
          7111 => x"5c",
          7112 => x"54",
          7113 => x"8e",
          7114 => x"07",
          7115 => x"83",
          7116 => x"58",
          7117 => x"18",
          7118 => x"75",
          7119 => x"18",
          7120 => x"39",
          7121 => x"54",
          7122 => x"2e",
          7123 => x"86",
          7124 => x"a0",
          7125 => x"88",
          7126 => x"06",
          7127 => x"82",
          7128 => x"06",
          7129 => x"06",
          7130 => x"2e",
          7131 => x"83",
          7132 => x"83",
          7133 => x"06",
          7134 => x"82",
          7135 => x"81",
          7136 => x"06",
          7137 => x"9f",
          7138 => x"06",
          7139 => x"2e",
          7140 => x"90",
          7141 => x"82",
          7142 => x"06",
          7143 => x"80",
          7144 => x"76",
          7145 => x"76",
          7146 => x"7d",
          7147 => x"3f",
          7148 => x"08",
          7149 => x"56",
          7150 => x"d8",
          7151 => x"be",
          7152 => x"d8",
          7153 => x"09",
          7154 => x"e8",
          7155 => x"2a",
          7156 => x"76",
          7157 => x"51",
          7158 => x"2e",
          7159 => x"81",
          7160 => x"80",
          7161 => x"38",
          7162 => x"ab",
          7163 => x"56",
          7164 => x"74",
          7165 => x"73",
          7166 => x"56",
          7167 => x"82",
          7168 => x"06",
          7169 => x"ac",
          7170 => x"33",
          7171 => x"70",
          7172 => x"55",
          7173 => x"2e",
          7174 => x"1e",
          7175 => x"06",
          7176 => x"05",
          7177 => x"e4",
          7178 => x"d6",
          7179 => x"1f",
          7180 => x"39",
          7181 => x"d8",
          7182 => x"0d",
          7183 => x"0d",
          7184 => x"7b",
          7185 => x"73",
          7186 => x"55",
          7187 => x"2e",
          7188 => x"75",
          7189 => x"57",
          7190 => x"26",
          7191 => x"ba",
          7192 => x"70",
          7193 => x"ba",
          7194 => x"06",
          7195 => x"73",
          7196 => x"70",
          7197 => x"51",
          7198 => x"89",
          7199 => x"82",
          7200 => x"ff",
          7201 => x"56",
          7202 => x"2e",
          7203 => x"80",
          7204 => x"c4",
          7205 => x"08",
          7206 => x"76",
          7207 => x"58",
          7208 => x"81",
          7209 => x"ff",
          7210 => x"53",
          7211 => x"26",
          7212 => x"13",
          7213 => x"06",
          7214 => x"9f",
          7215 => x"99",
          7216 => x"e0",
          7217 => x"ff",
          7218 => x"72",
          7219 => x"2a",
          7220 => x"72",
          7221 => x"06",
          7222 => x"ff",
          7223 => x"30",
          7224 => x"70",
          7225 => x"07",
          7226 => x"9f",
          7227 => x"54",
          7228 => x"80",
          7229 => x"81",
          7230 => x"59",
          7231 => x"25",
          7232 => x"8b",
          7233 => x"24",
          7234 => x"76",
          7235 => x"78",
          7236 => x"82",
          7237 => x"51",
          7238 => x"d8",
          7239 => x"0d",
          7240 => x"0d",
          7241 => x"0b",
          7242 => x"ff",
          7243 => x"0c",
          7244 => x"51",
          7245 => x"84",
          7246 => x"d8",
          7247 => x"38",
          7248 => x"51",
          7249 => x"82",
          7250 => x"83",
          7251 => x"54",
          7252 => x"82",
          7253 => x"09",
          7254 => x"e3",
          7255 => x"b8",
          7256 => x"57",
          7257 => x"2e",
          7258 => x"83",
          7259 => x"74",
          7260 => x"70",
          7261 => x"25",
          7262 => x"51",
          7263 => x"38",
          7264 => x"2e",
          7265 => x"b5",
          7266 => x"82",
          7267 => x"80",
          7268 => x"cf",
          7269 => x"d6",
          7270 => x"82",
          7271 => x"80",
          7272 => x"85",
          7273 => x"88",
          7274 => x"16",
          7275 => x"3f",
          7276 => x"08",
          7277 => x"d8",
          7278 => x"83",
          7279 => x"74",
          7280 => x"0c",
          7281 => x"04",
          7282 => x"61",
          7283 => x"80",
          7284 => x"58",
          7285 => x"0c",
          7286 => x"e1",
          7287 => x"d8",
          7288 => x"56",
          7289 => x"d6",
          7290 => x"87",
          7291 => x"d6",
          7292 => x"29",
          7293 => x"05",
          7294 => x"53",
          7295 => x"80",
          7296 => x"38",
          7297 => x"76",
          7298 => x"74",
          7299 => x"72",
          7300 => x"38",
          7301 => x"51",
          7302 => x"82",
          7303 => x"81",
          7304 => x"81",
          7305 => x"72",
          7306 => x"80",
          7307 => x"38",
          7308 => x"70",
          7309 => x"53",
          7310 => x"86",
          7311 => x"af",
          7312 => x"34",
          7313 => x"34",
          7314 => x"14",
          7315 => x"88",
          7316 => x"d8",
          7317 => x"06",
          7318 => x"54",
          7319 => x"72",
          7320 => x"76",
          7321 => x"38",
          7322 => x"70",
          7323 => x"53",
          7324 => x"85",
          7325 => x"70",
          7326 => x"5b",
          7327 => x"82",
          7328 => x"81",
          7329 => x"76",
          7330 => x"81",
          7331 => x"38",
          7332 => x"56",
          7333 => x"83",
          7334 => x"70",
          7335 => x"80",
          7336 => x"83",
          7337 => x"cb",
          7338 => x"d6",
          7339 => x"76",
          7340 => x"05",
          7341 => x"16",
          7342 => x"56",
          7343 => x"d7",
          7344 => x"8d",
          7345 => x"72",
          7346 => x"54",
          7347 => x"57",
          7348 => x"95",
          7349 => x"73",
          7350 => x"3f",
          7351 => x"08",
          7352 => x"57",
          7353 => x"89",
          7354 => x"56",
          7355 => x"d7",
          7356 => x"76",
          7357 => x"f9",
          7358 => x"76",
          7359 => x"f1",
          7360 => x"14",
          7361 => x"3f",
          7362 => x"08",
          7363 => x"06",
          7364 => x"80",
          7365 => x"06",
          7366 => x"80",
          7367 => x"ca",
          7368 => x"d6",
          7369 => x"ff",
          7370 => x"77",
          7371 => x"dc",
          7372 => x"b3",
          7373 => x"d8",
          7374 => x"a0",
          7375 => x"c8",
          7376 => x"15",
          7377 => x"14",
          7378 => x"70",
          7379 => x"51",
          7380 => x"56",
          7381 => x"84",
          7382 => x"81",
          7383 => x"71",
          7384 => x"16",
          7385 => x"53",
          7386 => x"23",
          7387 => x"8b",
          7388 => x"73",
          7389 => x"80",
          7390 => x"8d",
          7391 => x"39",
          7392 => x"51",
          7393 => x"82",
          7394 => x"53",
          7395 => x"08",
          7396 => x"72",
          7397 => x"8d",
          7398 => x"d5",
          7399 => x"14",
          7400 => x"3f",
          7401 => x"08",
          7402 => x"06",
          7403 => x"38",
          7404 => x"51",
          7405 => x"82",
          7406 => x"55",
          7407 => x"51",
          7408 => x"82",
          7409 => x"83",
          7410 => x"53",
          7411 => x"80",
          7412 => x"38",
          7413 => x"78",
          7414 => x"2a",
          7415 => x"78",
          7416 => x"8d",
          7417 => x"22",
          7418 => x"31",
          7419 => x"c1",
          7420 => x"d8",
          7421 => x"d6",
          7422 => x"2e",
          7423 => x"82",
          7424 => x"80",
          7425 => x"f5",
          7426 => x"83",
          7427 => x"ff",
          7428 => x"38",
          7429 => x"9f",
          7430 => x"38",
          7431 => x"39",
          7432 => x"80",
          7433 => x"38",
          7434 => x"9c",
          7435 => x"a4",
          7436 => x"1c",
          7437 => x"0c",
          7438 => x"17",
          7439 => x"76",
          7440 => x"81",
          7441 => x"80",
          7442 => x"c8",
          7443 => x"d6",
          7444 => x"ff",
          7445 => x"8d",
          7446 => x"95",
          7447 => x"91",
          7448 => x"14",
          7449 => x"3f",
          7450 => x"08",
          7451 => x"74",
          7452 => x"a2",
          7453 => x"79",
          7454 => x"f5",
          7455 => x"ac",
          7456 => x"15",
          7457 => x"2e",
          7458 => x"10",
          7459 => x"2a",
          7460 => x"05",
          7461 => x"ff",
          7462 => x"53",
          7463 => x"a0",
          7464 => x"81",
          7465 => x"0b",
          7466 => x"ff",
          7467 => x"0c",
          7468 => x"84",
          7469 => x"83",
          7470 => x"06",
          7471 => x"80",
          7472 => x"c7",
          7473 => x"d6",
          7474 => x"ff",
          7475 => x"72",
          7476 => x"81",
          7477 => x"38",
          7478 => x"73",
          7479 => x"3f",
          7480 => x"08",
          7481 => x"82",
          7482 => x"84",
          7483 => x"b6",
          7484 => x"dc",
          7485 => x"d8",
          7486 => x"ff",
          7487 => x"82",
          7488 => x"09",
          7489 => x"c8",
          7490 => x"51",
          7491 => x"82",
          7492 => x"84",
          7493 => x"d2",
          7494 => x"06",
          7495 => x"9c",
          7496 => x"c3",
          7497 => x"d8",
          7498 => x"85",
          7499 => x"09",
          7500 => x"38",
          7501 => x"51",
          7502 => x"82",
          7503 => x"94",
          7504 => x"a4",
          7505 => x"9f",
          7506 => x"d8",
          7507 => x"0c",
          7508 => x"82",
          7509 => x"81",
          7510 => x"82",
          7511 => x"72",
          7512 => x"82",
          7513 => x"8c",
          7514 => x"0b",
          7515 => x"80",
          7516 => x"d6",
          7517 => x"3d",
          7518 => x"3d",
          7519 => x"89",
          7520 => x"2e",
          7521 => x"08",
          7522 => x"2e",
          7523 => x"33",
          7524 => x"2e",
          7525 => x"13",
          7526 => x"22",
          7527 => x"76",
          7528 => x"06",
          7529 => x"13",
          7530 => x"bf",
          7531 => x"d6",
          7532 => x"06",
          7533 => x"38",
          7534 => x"54",
          7535 => x"80",
          7536 => x"71",
          7537 => x"82",
          7538 => x"87",
          7539 => x"fa",
          7540 => x"ab",
          7541 => x"58",
          7542 => x"05",
          7543 => x"dd",
          7544 => x"80",
          7545 => x"d8",
          7546 => x"38",
          7547 => x"08",
          7548 => x"ee",
          7549 => x"08",
          7550 => x"80",
          7551 => x"80",
          7552 => x"54",
          7553 => x"84",
          7554 => x"34",
          7555 => x"75",
          7556 => x"2e",
          7557 => x"53",
          7558 => x"53",
          7559 => x"f7",
          7560 => x"d6",
          7561 => x"73",
          7562 => x"0c",
          7563 => x"04",
          7564 => x"68",
          7565 => x"80",
          7566 => x"59",
          7567 => x"78",
          7568 => x"c8",
          7569 => x"06",
          7570 => x"3d",
          7571 => x"9a",
          7572 => x"52",
          7573 => x"3f",
          7574 => x"08",
          7575 => x"d8",
          7576 => x"38",
          7577 => x"52",
          7578 => x"52",
          7579 => x"3f",
          7580 => x"08",
          7581 => x"d8",
          7582 => x"02",
          7583 => x"33",
          7584 => x"55",
          7585 => x"25",
          7586 => x"55",
          7587 => x"54",
          7588 => x"81",
          7589 => x"80",
          7590 => x"74",
          7591 => x"81",
          7592 => x"75",
          7593 => x"3f",
          7594 => x"08",
          7595 => x"02",
          7596 => x"91",
          7597 => x"81",
          7598 => x"82",
          7599 => x"06",
          7600 => x"80",
          7601 => x"88",
          7602 => x"39",
          7603 => x"58",
          7604 => x"38",
          7605 => x"70",
          7606 => x"54",
          7607 => x"81",
          7608 => x"52",
          7609 => x"b0",
          7610 => x"d8",
          7611 => x"88",
          7612 => x"62",
          7613 => x"c3",
          7614 => x"54",
          7615 => x"15",
          7616 => x"62",
          7617 => x"d7",
          7618 => x"52",
          7619 => x"51",
          7620 => x"7a",
          7621 => x"83",
          7622 => x"80",
          7623 => x"38",
          7624 => x"08",
          7625 => x"53",
          7626 => x"3d",
          7627 => x"cc",
          7628 => x"d6",
          7629 => x"82",
          7630 => x"82",
          7631 => x"39",
          7632 => x"38",
          7633 => x"33",
          7634 => x"70",
          7635 => x"55",
          7636 => x"2e",
          7637 => x"55",
          7638 => x"77",
          7639 => x"81",
          7640 => x"73",
          7641 => x"38",
          7642 => x"54",
          7643 => x"a0",
          7644 => x"82",
          7645 => x"52",
          7646 => x"ae",
          7647 => x"d8",
          7648 => x"18",
          7649 => x"55",
          7650 => x"d8",
          7651 => x"38",
          7652 => x"70",
          7653 => x"54",
          7654 => x"86",
          7655 => x"c0",
          7656 => x"b4",
          7657 => x"1b",
          7658 => x"1b",
          7659 => x"70",
          7660 => x"e4",
          7661 => x"d8",
          7662 => x"d8",
          7663 => x"0c",
          7664 => x"52",
          7665 => x"3f",
          7666 => x"08",
          7667 => x"08",
          7668 => x"77",
          7669 => x"86",
          7670 => x"1a",
          7671 => x"1a",
          7672 => x"91",
          7673 => x"0b",
          7674 => x"80",
          7675 => x"0c",
          7676 => x"70",
          7677 => x"54",
          7678 => x"81",
          7679 => x"d6",
          7680 => x"2e",
          7681 => x"82",
          7682 => x"94",
          7683 => x"17",
          7684 => x"2b",
          7685 => x"57",
          7686 => x"52",
          7687 => x"aa",
          7688 => x"d8",
          7689 => x"d6",
          7690 => x"26",
          7691 => x"55",
          7692 => x"08",
          7693 => x"81",
          7694 => x"79",
          7695 => x"31",
          7696 => x"70",
          7697 => x"25",
          7698 => x"76",
          7699 => x"81",
          7700 => x"55",
          7701 => x"38",
          7702 => x"0c",
          7703 => x"75",
          7704 => x"54",
          7705 => x"a2",
          7706 => x"7a",
          7707 => x"3f",
          7708 => x"08",
          7709 => x"55",
          7710 => x"89",
          7711 => x"d8",
          7712 => x"1a",
          7713 => x"80",
          7714 => x"54",
          7715 => x"d8",
          7716 => x"0d",
          7717 => x"0d",
          7718 => x"64",
          7719 => x"59",
          7720 => x"90",
          7721 => x"52",
          7722 => x"ce",
          7723 => x"d8",
          7724 => x"d6",
          7725 => x"38",
          7726 => x"55",
          7727 => x"86",
          7728 => x"82",
          7729 => x"19",
          7730 => x"55",
          7731 => x"80",
          7732 => x"38",
          7733 => x"0b",
          7734 => x"82",
          7735 => x"39",
          7736 => x"1a",
          7737 => x"82",
          7738 => x"19",
          7739 => x"08",
          7740 => x"7c",
          7741 => x"74",
          7742 => x"2e",
          7743 => x"94",
          7744 => x"83",
          7745 => x"56",
          7746 => x"38",
          7747 => x"22",
          7748 => x"89",
          7749 => x"55",
          7750 => x"75",
          7751 => x"19",
          7752 => x"39",
          7753 => x"52",
          7754 => x"9e",
          7755 => x"d8",
          7756 => x"75",
          7757 => x"38",
          7758 => x"ff",
          7759 => x"98",
          7760 => x"19",
          7761 => x"51",
          7762 => x"82",
          7763 => x"80",
          7764 => x"38",
          7765 => x"08",
          7766 => x"2a",
          7767 => x"80",
          7768 => x"38",
          7769 => x"8a",
          7770 => x"5c",
          7771 => x"27",
          7772 => x"7a",
          7773 => x"54",
          7774 => x"52",
          7775 => x"51",
          7776 => x"3f",
          7777 => x"08",
          7778 => x"7e",
          7779 => x"56",
          7780 => x"2e",
          7781 => x"16",
          7782 => x"55",
          7783 => x"95",
          7784 => x"53",
          7785 => x"b4",
          7786 => x"31",
          7787 => x"05",
          7788 => x"ab",
          7789 => x"2b",
          7790 => x"76",
          7791 => x"94",
          7792 => x"ff",
          7793 => x"71",
          7794 => x"7b",
          7795 => x"38",
          7796 => x"19",
          7797 => x"51",
          7798 => x"82",
          7799 => x"fd",
          7800 => x"53",
          7801 => x"83",
          7802 => x"b8",
          7803 => x"51",
          7804 => x"3f",
          7805 => x"7e",
          7806 => x"0c",
          7807 => x"1b",
          7808 => x"1c",
          7809 => x"fd",
          7810 => x"56",
          7811 => x"d8",
          7812 => x"0d",
          7813 => x"0d",
          7814 => x"64",
          7815 => x"58",
          7816 => x"90",
          7817 => x"52",
          7818 => x"ce",
          7819 => x"d8",
          7820 => x"d6",
          7821 => x"38",
          7822 => x"55",
          7823 => x"86",
          7824 => x"83",
          7825 => x"18",
          7826 => x"2a",
          7827 => x"51",
          7828 => x"56",
          7829 => x"83",
          7830 => x"39",
          7831 => x"19",
          7832 => x"83",
          7833 => x"0b",
          7834 => x"81",
          7835 => x"39",
          7836 => x"7c",
          7837 => x"74",
          7838 => x"38",
          7839 => x"7b",
          7840 => x"f2",
          7841 => x"08",
          7842 => x"06",
          7843 => x"82",
          7844 => x"8a",
          7845 => x"05",
          7846 => x"06",
          7847 => x"bf",
          7848 => x"38",
          7849 => x"55",
          7850 => x"7a",
          7851 => x"98",
          7852 => x"77",
          7853 => x"3f",
          7854 => x"08",
          7855 => x"d8",
          7856 => x"82",
          7857 => x"81",
          7858 => x"38",
          7859 => x"ff",
          7860 => x"98",
          7861 => x"18",
          7862 => x"74",
          7863 => x"7e",
          7864 => x"08",
          7865 => x"2e",
          7866 => x"8e",
          7867 => x"ff",
          7868 => x"82",
          7869 => x"fe",
          7870 => x"18",
          7871 => x"51",
          7872 => x"82",
          7873 => x"80",
          7874 => x"38",
          7875 => x"08",
          7876 => x"2a",
          7877 => x"80",
          7878 => x"38",
          7879 => x"8a",
          7880 => x"5b",
          7881 => x"27",
          7882 => x"7b",
          7883 => x"54",
          7884 => x"52",
          7885 => x"51",
          7886 => x"3f",
          7887 => x"08",
          7888 => x"7e",
          7889 => x"78",
          7890 => x"74",
          7891 => x"38",
          7892 => x"b4",
          7893 => x"31",
          7894 => x"05",
          7895 => x"51",
          7896 => x"3f",
          7897 => x"0b",
          7898 => x"78",
          7899 => x"80",
          7900 => x"18",
          7901 => x"08",
          7902 => x"7e",
          7903 => x"ba",
          7904 => x"d8",
          7905 => x"38",
          7906 => x"12",
          7907 => x"9c",
          7908 => x"18",
          7909 => x"06",
          7910 => x"31",
          7911 => x"76",
          7912 => x"7b",
          7913 => x"08",
          7914 => x"ff",
          7915 => x"82",
          7916 => x"fd",
          7917 => x"53",
          7918 => x"18",
          7919 => x"06",
          7920 => x"51",
          7921 => x"3f",
          7922 => x"0b",
          7923 => x"7b",
          7924 => x"08",
          7925 => x"76",
          7926 => x"08",
          7927 => x"1c",
          7928 => x"08",
          7929 => x"5c",
          7930 => x"83",
          7931 => x"74",
          7932 => x"fd",
          7933 => x"18",
          7934 => x"07",
          7935 => x"19",
          7936 => x"75",
          7937 => x"0c",
          7938 => x"04",
          7939 => x"7a",
          7940 => x"05",
          7941 => x"56",
          7942 => x"82",
          7943 => x"57",
          7944 => x"08",
          7945 => x"90",
          7946 => x"86",
          7947 => x"06",
          7948 => x"73",
          7949 => x"ee",
          7950 => x"08",
          7951 => x"ff",
          7952 => x"82",
          7953 => x"57",
          7954 => x"08",
          7955 => x"a4",
          7956 => x"11",
          7957 => x"55",
          7958 => x"16",
          7959 => x"08",
          7960 => x"75",
          7961 => x"e9",
          7962 => x"08",
          7963 => x"51",
          7964 => x"3f",
          7965 => x"0a",
          7966 => x"51",
          7967 => x"3f",
          7968 => x"15",
          7969 => x"8a",
          7970 => x"81",
          7971 => x"34",
          7972 => x"bb",
          7973 => x"d6",
          7974 => x"17",
          7975 => x"06",
          7976 => x"90",
          7977 => x"82",
          7978 => x"8a",
          7979 => x"fc",
          7980 => x"70",
          7981 => x"d4",
          7982 => x"d8",
          7983 => x"d6",
          7984 => x"38",
          7985 => x"05",
          7986 => x"f1",
          7987 => x"d6",
          7988 => x"82",
          7989 => x"87",
          7990 => x"d8",
          7991 => x"72",
          7992 => x"0c",
          7993 => x"04",
          7994 => x"84",
          7995 => x"cd",
          7996 => x"80",
          7997 => x"d8",
          7998 => x"38",
          7999 => x"08",
          8000 => x"34",
          8001 => x"82",
          8002 => x"83",
          8003 => x"ee",
          8004 => x"53",
          8005 => x"05",
          8006 => x"51",
          8007 => x"82",
          8008 => x"55",
          8009 => x"08",
          8010 => x"76",
          8011 => x"94",
          8012 => x"51",
          8013 => x"82",
          8014 => x"55",
          8015 => x"08",
          8016 => x"80",
          8017 => x"70",
          8018 => x"56",
          8019 => x"89",
          8020 => x"98",
          8021 => x"b2",
          8022 => x"05",
          8023 => x"2a",
          8024 => x"51",
          8025 => x"80",
          8026 => x"76",
          8027 => x"52",
          8028 => x"3f",
          8029 => x"08",
          8030 => x"8e",
          8031 => x"d8",
          8032 => x"09",
          8033 => x"38",
          8034 => x"82",
          8035 => x"94",
          8036 => x"ff",
          8037 => x"80",
          8038 => x"80",
          8039 => x"5b",
          8040 => x"34",
          8041 => x"df",
          8042 => x"05",
          8043 => x"3d",
          8044 => x"3f",
          8045 => x"08",
          8046 => x"d8",
          8047 => x"38",
          8048 => x"3d",
          8049 => x"98",
          8050 => x"d8",
          8051 => x"58",
          8052 => x"08",
          8053 => x"2e",
          8054 => x"a0",
          8055 => x"3d",
          8056 => x"c4",
          8057 => x"d6",
          8058 => x"82",
          8059 => x"82",
          8060 => x"d9",
          8061 => x"7b",
          8062 => x"ae",
          8063 => x"d8",
          8064 => x"d6",
          8065 => x"d8",
          8066 => x"3d",
          8067 => x"51",
          8068 => x"82",
          8069 => x"80",
          8070 => x"76",
          8071 => x"c4",
          8072 => x"d6",
          8073 => x"82",
          8074 => x"82",
          8075 => x"52",
          8076 => x"fa",
          8077 => x"d8",
          8078 => x"d6",
          8079 => x"38",
          8080 => x"08",
          8081 => x"c8",
          8082 => x"82",
          8083 => x"2e",
          8084 => x"52",
          8085 => x"ac",
          8086 => x"d8",
          8087 => x"d6",
          8088 => x"2e",
          8089 => x"84",
          8090 => x"06",
          8091 => x"57",
          8092 => x"76",
          8093 => x"80",
          8094 => x"b8",
          8095 => x"51",
          8096 => x"76",
          8097 => x"11",
          8098 => x"51",
          8099 => x"73",
          8100 => x"38",
          8101 => x"05",
          8102 => x"81",
          8103 => x"56",
          8104 => x"f5",
          8105 => x"54",
          8106 => x"81",
          8107 => x"80",
          8108 => x"78",
          8109 => x"55",
          8110 => x"e1",
          8111 => x"ff",
          8112 => x"58",
          8113 => x"74",
          8114 => x"75",
          8115 => x"18",
          8116 => x"08",
          8117 => x"af",
          8118 => x"f4",
          8119 => x"2e",
          8120 => x"8d",
          8121 => x"80",
          8122 => x"11",
          8123 => x"74",
          8124 => x"82",
          8125 => x"70",
          8126 => x"c7",
          8127 => x"08",
          8128 => x"5c",
          8129 => x"73",
          8130 => x"38",
          8131 => x"1a",
          8132 => x"55",
          8133 => x"38",
          8134 => x"73",
          8135 => x"38",
          8136 => x"76",
          8137 => x"74",
          8138 => x"33",
          8139 => x"05",
          8140 => x"15",
          8141 => x"ba",
          8142 => x"05",
          8143 => x"ff",
          8144 => x"06",
          8145 => x"57",
          8146 => x"e0",
          8147 => x"81",
          8148 => x"73",
          8149 => x"81",
          8150 => x"7a",
          8151 => x"38",
          8152 => x"76",
          8153 => x"0c",
          8154 => x"0d",
          8155 => x"0d",
          8156 => x"3d",
          8157 => x"71",
          8158 => x"eb",
          8159 => x"d6",
          8160 => x"82",
          8161 => x"82",
          8162 => x"15",
          8163 => x"82",
          8164 => x"15",
          8165 => x"76",
          8166 => x"90",
          8167 => x"81",
          8168 => x"06",
          8169 => x"72",
          8170 => x"56",
          8171 => x"54",
          8172 => x"17",
          8173 => x"78",
          8174 => x"38",
          8175 => x"22",
          8176 => x"59",
          8177 => x"78",
          8178 => x"76",
          8179 => x"51",
          8180 => x"3f",
          8181 => x"08",
          8182 => x"54",
          8183 => x"53",
          8184 => x"3f",
          8185 => x"08",
          8186 => x"38",
          8187 => x"75",
          8188 => x"18",
          8189 => x"31",
          8190 => x"57",
          8191 => x"b2",
          8192 => x"08",
          8193 => x"38",
          8194 => x"51",
          8195 => x"3f",
          8196 => x"08",
          8197 => x"d8",
          8198 => x"81",
          8199 => x"d6",
          8200 => x"2e",
          8201 => x"82",
          8202 => x"88",
          8203 => x"98",
          8204 => x"80",
          8205 => x"38",
          8206 => x"80",
          8207 => x"77",
          8208 => x"08",
          8209 => x"0c",
          8210 => x"70",
          8211 => x"81",
          8212 => x"5a",
          8213 => x"2e",
          8214 => x"52",
          8215 => x"bb",
          8216 => x"d6",
          8217 => x"82",
          8218 => x"95",
          8219 => x"d8",
          8220 => x"39",
          8221 => x"51",
          8222 => x"3f",
          8223 => x"08",
          8224 => x"2e",
          8225 => x"74",
          8226 => x"79",
          8227 => x"14",
          8228 => x"38",
          8229 => x"0c",
          8230 => x"94",
          8231 => x"94",
          8232 => x"83",
          8233 => x"72",
          8234 => x"38",
          8235 => x"51",
          8236 => x"3f",
          8237 => x"08",
          8238 => x"0b",
          8239 => x"82",
          8240 => x"39",
          8241 => x"16",
          8242 => x"bb",
          8243 => x"2a",
          8244 => x"08",
          8245 => x"15",
          8246 => x"15",
          8247 => x"90",
          8248 => x"16",
          8249 => x"33",
          8250 => x"53",
          8251 => x"34",
          8252 => x"06",
          8253 => x"2e",
          8254 => x"9c",
          8255 => x"85",
          8256 => x"16",
          8257 => x"72",
          8258 => x"0c",
          8259 => x"04",
          8260 => x"79",
          8261 => x"75",
          8262 => x"8b",
          8263 => x"89",
          8264 => x"52",
          8265 => x"05",
          8266 => x"3f",
          8267 => x"08",
          8268 => x"d8",
          8269 => x"38",
          8270 => x"7a",
          8271 => x"d5",
          8272 => x"d6",
          8273 => x"82",
          8274 => x"80",
          8275 => x"16",
          8276 => x"2b",
          8277 => x"74",
          8278 => x"86",
          8279 => x"84",
          8280 => x"06",
          8281 => x"73",
          8282 => x"38",
          8283 => x"52",
          8284 => x"a4",
          8285 => x"d8",
          8286 => x"0c",
          8287 => x"14",
          8288 => x"23",
          8289 => x"51",
          8290 => x"3f",
          8291 => x"08",
          8292 => x"2e",
          8293 => x"85",
          8294 => x"86",
          8295 => x"2e",
          8296 => x"76",
          8297 => x"73",
          8298 => x"0c",
          8299 => x"04",
          8300 => x"76",
          8301 => x"05",
          8302 => x"53",
          8303 => x"82",
          8304 => x"87",
          8305 => x"d8",
          8306 => x"86",
          8307 => x"fb",
          8308 => x"79",
          8309 => x"05",
          8310 => x"56",
          8311 => x"3f",
          8312 => x"08",
          8313 => x"d8",
          8314 => x"38",
          8315 => x"82",
          8316 => x"52",
          8317 => x"bc",
          8318 => x"d6",
          8319 => x"80",
          8320 => x"d6",
          8321 => x"73",
          8322 => x"3f",
          8323 => x"08",
          8324 => x"d8",
          8325 => x"09",
          8326 => x"38",
          8327 => x"39",
          8328 => x"08",
          8329 => x"52",
          8330 => x"ba",
          8331 => x"73",
          8332 => x"d0",
          8333 => x"d8",
          8334 => x"70",
          8335 => x"07",
          8336 => x"82",
          8337 => x"06",
          8338 => x"54",
          8339 => x"d8",
          8340 => x"0d",
          8341 => x"0d",
          8342 => x"53",
          8343 => x"53",
          8344 => x"56",
          8345 => x"82",
          8346 => x"55",
          8347 => x"08",
          8348 => x"52",
          8349 => x"ea",
          8350 => x"d8",
          8351 => x"d6",
          8352 => x"38",
          8353 => x"05",
          8354 => x"2b",
          8355 => x"80",
          8356 => x"86",
          8357 => x"76",
          8358 => x"38",
          8359 => x"51",
          8360 => x"74",
          8361 => x"0c",
          8362 => x"04",
          8363 => x"63",
          8364 => x"80",
          8365 => x"ec",
          8366 => x"3d",
          8367 => x"3f",
          8368 => x"08",
          8369 => x"d8",
          8370 => x"38",
          8371 => x"73",
          8372 => x"08",
          8373 => x"13",
          8374 => x"58",
          8375 => x"26",
          8376 => x"7c",
          8377 => x"39",
          8378 => x"ce",
          8379 => x"81",
          8380 => x"d6",
          8381 => x"33",
          8382 => x"81",
          8383 => x"06",
          8384 => x"82",
          8385 => x"76",
          8386 => x"f0",
          8387 => x"b0",
          8388 => x"d6",
          8389 => x"2e",
          8390 => x"d6",
          8391 => x"2e",
          8392 => x"d6",
          8393 => x"70",
          8394 => x"08",
          8395 => x"7a",
          8396 => x"7f",
          8397 => x"54",
          8398 => x"77",
          8399 => x"80",
          8400 => x"15",
          8401 => x"d8",
          8402 => x"75",
          8403 => x"52",
          8404 => x"52",
          8405 => x"d2",
          8406 => x"d8",
          8407 => x"d6",
          8408 => x"d6",
          8409 => x"33",
          8410 => x"1a",
          8411 => x"54",
          8412 => x"09",
          8413 => x"38",
          8414 => x"ff",
          8415 => x"82",
          8416 => x"83",
          8417 => x"70",
          8418 => x"25",
          8419 => x"59",
          8420 => x"9b",
          8421 => x"51",
          8422 => x"3f",
          8423 => x"08",
          8424 => x"70",
          8425 => x"25",
          8426 => x"59",
          8427 => x"75",
          8428 => x"7a",
          8429 => x"ff",
          8430 => x"7c",
          8431 => x"94",
          8432 => x"11",
          8433 => x"56",
          8434 => x"15",
          8435 => x"d6",
          8436 => x"3d",
          8437 => x"3d",
          8438 => x"3d",
          8439 => x"70",
          8440 => x"96",
          8441 => x"d8",
          8442 => x"d6",
          8443 => x"aa",
          8444 => x"33",
          8445 => x"a2",
          8446 => x"33",
          8447 => x"70",
          8448 => x"55",
          8449 => x"73",
          8450 => x"90",
          8451 => x"08",
          8452 => x"18",
          8453 => x"82",
          8454 => x"38",
          8455 => x"08",
          8456 => x"08",
          8457 => x"ff",
          8458 => x"82",
          8459 => x"74",
          8460 => x"56",
          8461 => x"98",
          8462 => x"76",
          8463 => x"8a",
          8464 => x"d8",
          8465 => x"09",
          8466 => x"38",
          8467 => x"d6",
          8468 => x"2e",
          8469 => x"85",
          8470 => x"a4",
          8471 => x"38",
          8472 => x"d6",
          8473 => x"15",
          8474 => x"38",
          8475 => x"53",
          8476 => x"08",
          8477 => x"ff",
          8478 => x"82",
          8479 => x"56",
          8480 => x"8c",
          8481 => x"17",
          8482 => x"07",
          8483 => x"18",
          8484 => x"2e",
          8485 => x"91",
          8486 => x"55",
          8487 => x"d8",
          8488 => x"0d",
          8489 => x"0d",
          8490 => x"3d",
          8491 => x"52",
          8492 => x"da",
          8493 => x"d6",
          8494 => x"82",
          8495 => x"81",
          8496 => x"46",
          8497 => x"52",
          8498 => x"52",
          8499 => x"3f",
          8500 => x"08",
          8501 => x"d8",
          8502 => x"38",
          8503 => x"05",
          8504 => x"2a",
          8505 => x"51",
          8506 => x"55",
          8507 => x"38",
          8508 => x"54",
          8509 => x"81",
          8510 => x"80",
          8511 => x"70",
          8512 => x"54",
          8513 => x"81",
          8514 => x"52",
          8515 => x"bb",
          8516 => x"d6",
          8517 => x"84",
          8518 => x"06",
          8519 => x"73",
          8520 => x"d6",
          8521 => x"82",
          8522 => x"98",
          8523 => x"81",
          8524 => x"5a",
          8525 => x"08",
          8526 => x"8a",
          8527 => x"54",
          8528 => x"3f",
          8529 => x"08",
          8530 => x"d8",
          8531 => x"38",
          8532 => x"08",
          8533 => x"ff",
          8534 => x"82",
          8535 => x"55",
          8536 => x"08",
          8537 => x"55",
          8538 => x"82",
          8539 => x"84",
          8540 => x"82",
          8541 => x"80",
          8542 => x"51",
          8543 => x"82",
          8544 => x"82",
          8545 => x"30",
          8546 => x"d8",
          8547 => x"25",
          8548 => x"75",
          8549 => x"38",
          8550 => x"90",
          8551 => x"75",
          8552 => x"ff",
          8553 => x"82",
          8554 => x"55",
          8555 => x"78",
          8556 => x"bd",
          8557 => x"d8",
          8558 => x"82",
          8559 => x"a2",
          8560 => x"e8",
          8561 => x"53",
          8562 => x"bc",
          8563 => x"3d",
          8564 => x"3f",
          8565 => x"08",
          8566 => x"d8",
          8567 => x"38",
          8568 => x"52",
          8569 => x"52",
          8570 => x"3f",
          8571 => x"08",
          8572 => x"d8",
          8573 => x"88",
          8574 => x"39",
          8575 => x"08",
          8576 => x"81",
          8577 => x"38",
          8578 => x"05",
          8579 => x"2a",
          8580 => x"55",
          8581 => x"81",
          8582 => x"5a",
          8583 => x"3d",
          8584 => x"ff",
          8585 => x"82",
          8586 => x"75",
          8587 => x"d6",
          8588 => x"38",
          8589 => x"d6",
          8590 => x"2e",
          8591 => x"83",
          8592 => x"82",
          8593 => x"ff",
          8594 => x"06",
          8595 => x"54",
          8596 => x"73",
          8597 => x"82",
          8598 => x"52",
          8599 => x"b2",
          8600 => x"d6",
          8601 => x"82",
          8602 => x"81",
          8603 => x"53",
          8604 => x"19",
          8605 => x"8a",
          8606 => x"ae",
          8607 => x"34",
          8608 => x"0b",
          8609 => x"34",
          8610 => x"0a",
          8611 => x"19",
          8612 => x"9c",
          8613 => x"78",
          8614 => x"51",
          8615 => x"3f",
          8616 => x"b8",
          8617 => x"d8",
          8618 => x"a4",
          8619 => x"54",
          8620 => x"d9",
          8621 => x"53",
          8622 => x"11",
          8623 => x"b8",
          8624 => x"54",
          8625 => x"15",
          8626 => x"ff",
          8627 => x"82",
          8628 => x"54",
          8629 => x"08",
          8630 => x"88",
          8631 => x"64",
          8632 => x"ff",
          8633 => x"75",
          8634 => x"78",
          8635 => x"e1",
          8636 => x"90",
          8637 => x"34",
          8638 => x"0b",
          8639 => x"78",
          8640 => x"ed",
          8641 => x"d8",
          8642 => x"39",
          8643 => x"52",
          8644 => x"ac",
          8645 => x"82",
          8646 => x"9a",
          8647 => x"d8",
          8648 => x"3d",
          8649 => x"d2",
          8650 => x"53",
          8651 => x"fc",
          8652 => x"3d",
          8653 => x"3f",
          8654 => x"08",
          8655 => x"d8",
          8656 => x"38",
          8657 => x"3d",
          8658 => x"3d",
          8659 => x"c9",
          8660 => x"d6",
          8661 => x"82",
          8662 => x"82",
          8663 => x"81",
          8664 => x"81",
          8665 => x"86",
          8666 => x"af",
          8667 => x"a5",
          8668 => x"aa",
          8669 => x"05",
          8670 => x"e3",
          8671 => x"77",
          8672 => x"70",
          8673 => x"a2",
          8674 => x"3d",
          8675 => x"51",
          8676 => x"82",
          8677 => x"55",
          8678 => x"08",
          8679 => x"a1",
          8680 => x"09",
          8681 => x"38",
          8682 => x"08",
          8683 => x"88",
          8684 => x"39",
          8685 => x"08",
          8686 => x"81",
          8687 => x"38",
          8688 => x"bd",
          8689 => x"d6",
          8690 => x"82",
          8691 => x"81",
          8692 => x"56",
          8693 => x"3d",
          8694 => x"52",
          8695 => x"ff",
          8696 => x"02",
          8697 => x"8b",
          8698 => x"16",
          8699 => x"2a",
          8700 => x"51",
          8701 => x"89",
          8702 => x"07",
          8703 => x"17",
          8704 => x"81",
          8705 => x"34",
          8706 => x"70",
          8707 => x"81",
          8708 => x"55",
          8709 => x"80",
          8710 => x"64",
          8711 => x"38",
          8712 => x"51",
          8713 => x"3f",
          8714 => x"08",
          8715 => x"ff",
          8716 => x"82",
          8717 => x"d8",
          8718 => x"80",
          8719 => x"d6",
          8720 => x"78",
          8721 => x"e2",
          8722 => x"d8",
          8723 => x"d8",
          8724 => x"55",
          8725 => x"08",
          8726 => x"81",
          8727 => x"73",
          8728 => x"81",
          8729 => x"63",
          8730 => x"76",
          8731 => x"e1",
          8732 => x"81",
          8733 => x"34",
          8734 => x"d6",
          8735 => x"38",
          8736 => x"e9",
          8737 => x"d8",
          8738 => x"d6",
          8739 => x"38",
          8740 => x"a3",
          8741 => x"d6",
          8742 => x"74",
          8743 => x"0c",
          8744 => x"04",
          8745 => x"02",
          8746 => x"33",
          8747 => x"80",
          8748 => x"57",
          8749 => x"96",
          8750 => x"52",
          8751 => x"d2",
          8752 => x"d6",
          8753 => x"82",
          8754 => x"80",
          8755 => x"5a",
          8756 => x"3d",
          8757 => x"c6",
          8758 => x"d6",
          8759 => x"82",
          8760 => x"b8",
          8761 => x"cf",
          8762 => x"a0",
          8763 => x"55",
          8764 => x"75",
          8765 => x"71",
          8766 => x"33",
          8767 => x"74",
          8768 => x"57",
          8769 => x"8b",
          8770 => x"54",
          8771 => x"15",
          8772 => x"ff",
          8773 => x"82",
          8774 => x"55",
          8775 => x"d8",
          8776 => x"0d",
          8777 => x"0d",
          8778 => x"53",
          8779 => x"05",
          8780 => x"51",
          8781 => x"82",
          8782 => x"55",
          8783 => x"08",
          8784 => x"76",
          8785 => x"94",
          8786 => x"51",
          8787 => x"82",
          8788 => x"55",
          8789 => x"08",
          8790 => x"80",
          8791 => x"81",
          8792 => x"86",
          8793 => x"38",
          8794 => x"86",
          8795 => x"90",
          8796 => x"54",
          8797 => x"ff",
          8798 => x"76",
          8799 => x"83",
          8800 => x"51",
          8801 => x"3f",
          8802 => x"08",
          8803 => x"d6",
          8804 => x"3d",
          8805 => x"3d",
          8806 => x"5c",
          8807 => x"99",
          8808 => x"52",
          8809 => x"d0",
          8810 => x"d6",
          8811 => x"d6",
          8812 => x"70",
          8813 => x"08",
          8814 => x"51",
          8815 => x"80",
          8816 => x"38",
          8817 => x"06",
          8818 => x"80",
          8819 => x"38",
          8820 => x"5f",
          8821 => x"3d",
          8822 => x"ff",
          8823 => x"82",
          8824 => x"57",
          8825 => x"08",
          8826 => x"74",
          8827 => x"ff",
          8828 => x"82",
          8829 => x"57",
          8830 => x"08",
          8831 => x"d6",
          8832 => x"d6",
          8833 => x"5b",
          8834 => x"18",
          8835 => x"18",
          8836 => x"74",
          8837 => x"81",
          8838 => x"78",
          8839 => x"8b",
          8840 => x"54",
          8841 => x"75",
          8842 => x"38",
          8843 => x"1b",
          8844 => x"55",
          8845 => x"2e",
          8846 => x"39",
          8847 => x"09",
          8848 => x"38",
          8849 => x"80",
          8850 => x"70",
          8851 => x"25",
          8852 => x"80",
          8853 => x"38",
          8854 => x"bc",
          8855 => x"11",
          8856 => x"ff",
          8857 => x"82",
          8858 => x"57",
          8859 => x"08",
          8860 => x"70",
          8861 => x"80",
          8862 => x"83",
          8863 => x"80",
          8864 => x"84",
          8865 => x"a7",
          8866 => x"b8",
          8867 => x"9b",
          8868 => x"d6",
          8869 => x"0c",
          8870 => x"d8",
          8871 => x"0d",
          8872 => x"0d",
          8873 => x"3d",
          8874 => x"52",
          8875 => x"ce",
          8876 => x"d6",
          8877 => x"d6",
          8878 => x"54",
          8879 => x"08",
          8880 => x"8b",
          8881 => x"8a",
          8882 => x"58",
          8883 => x"3f",
          8884 => x"33",
          8885 => x"9f",
          8886 => x"86",
          8887 => x"9d",
          8888 => x"9d",
          8889 => x"d6",
          8890 => x"ff",
          8891 => x"c4",
          8892 => x"d8",
          8893 => x"98",
          8894 => x"52",
          8895 => x"08",
          8896 => x"3f",
          8897 => x"08",
          8898 => x"06",
          8899 => x"2e",
          8900 => x"52",
          8901 => x"51",
          8902 => x"3f",
          8903 => x"08",
          8904 => x"ff",
          8905 => x"38",
          8906 => x"88",
          8907 => x"8a",
          8908 => x"38",
          8909 => x"e7",
          8910 => x"75",
          8911 => x"74",
          8912 => x"73",
          8913 => x"05",
          8914 => x"16",
          8915 => x"70",
          8916 => x"34",
          8917 => x"70",
          8918 => x"56",
          8919 => x"fe",
          8920 => x"3d",
          8921 => x"55",
          8922 => x"2e",
          8923 => x"75",
          8924 => x"38",
          8925 => x"55",
          8926 => x"33",
          8927 => x"a0",
          8928 => x"06",
          8929 => x"16",
          8930 => x"38",
          8931 => x"42",
          8932 => x"3d",
          8933 => x"ff",
          8934 => x"82",
          8935 => x"54",
          8936 => x"08",
          8937 => x"81",
          8938 => x"ff",
          8939 => x"82",
          8940 => x"54",
          8941 => x"08",
          8942 => x"80",
          8943 => x"54",
          8944 => x"80",
          8945 => x"d6",
          8946 => x"2e",
          8947 => x"80",
          8948 => x"54",
          8949 => x"80",
          8950 => x"52",
          8951 => x"ac",
          8952 => x"d6",
          8953 => x"82",
          8954 => x"b1",
          8955 => x"82",
          8956 => x"52",
          8957 => x"9a",
          8958 => x"54",
          8959 => x"15",
          8960 => x"77",
          8961 => x"ff",
          8962 => x"78",
          8963 => x"83",
          8964 => x"51",
          8965 => x"3f",
          8966 => x"08",
          8967 => x"74",
          8968 => x"0c",
          8969 => x"04",
          8970 => x"60",
          8971 => x"05",
          8972 => x"33",
          8973 => x"05",
          8974 => x"40",
          8975 => x"ba",
          8976 => x"d8",
          8977 => x"d6",
          8978 => x"bd",
          8979 => x"33",
          8980 => x"b5",
          8981 => x"2e",
          8982 => x"1a",
          8983 => x"90",
          8984 => x"33",
          8985 => x"70",
          8986 => x"55",
          8987 => x"38",
          8988 => x"97",
          8989 => x"82",
          8990 => x"58",
          8991 => x"7e",
          8992 => x"70",
          8993 => x"55",
          8994 => x"56",
          8995 => x"a1",
          8996 => x"7d",
          8997 => x"70",
          8998 => x"2a",
          8999 => x"08",
          9000 => x"08",
          9001 => x"5d",
          9002 => x"77",
          9003 => x"9c",
          9004 => x"26",
          9005 => x"57",
          9006 => x"59",
          9007 => x"52",
          9008 => x"9d",
          9009 => x"15",
          9010 => x"9c",
          9011 => x"26",
          9012 => x"55",
          9013 => x"08",
          9014 => x"99",
          9015 => x"d8",
          9016 => x"ff",
          9017 => x"d6",
          9018 => x"38",
          9019 => x"75",
          9020 => x"81",
          9021 => x"93",
          9022 => x"80",
          9023 => x"2e",
          9024 => x"ff",
          9025 => x"58",
          9026 => x"7d",
          9027 => x"38",
          9028 => x"55",
          9029 => x"b4",
          9030 => x"56",
          9031 => x"09",
          9032 => x"38",
          9033 => x"53",
          9034 => x"51",
          9035 => x"3f",
          9036 => x"08",
          9037 => x"d8",
          9038 => x"38",
          9039 => x"ff",
          9040 => x"5c",
          9041 => x"84",
          9042 => x"5c",
          9043 => x"12",
          9044 => x"80",
          9045 => x"78",
          9046 => x"7c",
          9047 => x"90",
          9048 => x"c0",
          9049 => x"90",
          9050 => x"15",
          9051 => x"94",
          9052 => x"54",
          9053 => x"91",
          9054 => x"31",
          9055 => x"84",
          9056 => x"07",
          9057 => x"16",
          9058 => x"73",
          9059 => x"0c",
          9060 => x"04",
          9061 => x"6b",
          9062 => x"05",
          9063 => x"33",
          9064 => x"5a",
          9065 => x"95",
          9066 => x"80",
          9067 => x"d8",
          9068 => x"f8",
          9069 => x"d8",
          9070 => x"82",
          9071 => x"70",
          9072 => x"74",
          9073 => x"38",
          9074 => x"82",
          9075 => x"81",
          9076 => x"81",
          9077 => x"ff",
          9078 => x"82",
          9079 => x"81",
          9080 => x"81",
          9081 => x"83",
          9082 => x"c0",
          9083 => x"2a",
          9084 => x"51",
          9085 => x"74",
          9086 => x"99",
          9087 => x"53",
          9088 => x"51",
          9089 => x"3f",
          9090 => x"08",
          9091 => x"55",
          9092 => x"92",
          9093 => x"80",
          9094 => x"38",
          9095 => x"06",
          9096 => x"2e",
          9097 => x"48",
          9098 => x"87",
          9099 => x"79",
          9100 => x"78",
          9101 => x"26",
          9102 => x"19",
          9103 => x"74",
          9104 => x"38",
          9105 => x"e4",
          9106 => x"2a",
          9107 => x"70",
          9108 => x"59",
          9109 => x"7a",
          9110 => x"56",
          9111 => x"80",
          9112 => x"51",
          9113 => x"74",
          9114 => x"99",
          9115 => x"53",
          9116 => x"51",
          9117 => x"3f",
          9118 => x"d6",
          9119 => x"ac",
          9120 => x"2a",
          9121 => x"82",
          9122 => x"43",
          9123 => x"83",
          9124 => x"66",
          9125 => x"60",
          9126 => x"90",
          9127 => x"31",
          9128 => x"80",
          9129 => x"8a",
          9130 => x"56",
          9131 => x"26",
          9132 => x"77",
          9133 => x"81",
          9134 => x"74",
          9135 => x"38",
          9136 => x"55",
          9137 => x"83",
          9138 => x"81",
          9139 => x"80",
          9140 => x"38",
          9141 => x"55",
          9142 => x"5e",
          9143 => x"89",
          9144 => x"5a",
          9145 => x"09",
          9146 => x"e1",
          9147 => x"38",
          9148 => x"57",
          9149 => x"c9",
          9150 => x"5a",
          9151 => x"9d",
          9152 => x"26",
          9153 => x"c9",
          9154 => x"10",
          9155 => x"22",
          9156 => x"74",
          9157 => x"38",
          9158 => x"ee",
          9159 => x"66",
          9160 => x"8d",
          9161 => x"d8",
          9162 => x"84",
          9163 => x"89",
          9164 => x"a0",
          9165 => x"82",
          9166 => x"fc",
          9167 => x"56",
          9168 => x"f0",
          9169 => x"80",
          9170 => x"d3",
          9171 => x"38",
          9172 => x"57",
          9173 => x"c8",
          9174 => x"5a",
          9175 => x"9d",
          9176 => x"26",
          9177 => x"c8",
          9178 => x"10",
          9179 => x"22",
          9180 => x"74",
          9181 => x"38",
          9182 => x"ee",
          9183 => x"66",
          9184 => x"ad",
          9185 => x"d8",
          9186 => x"05",
          9187 => x"d8",
          9188 => x"26",
          9189 => x"0b",
          9190 => x"08",
          9191 => x"d8",
          9192 => x"11",
          9193 => x"05",
          9194 => x"83",
          9195 => x"2a",
          9196 => x"a0",
          9197 => x"7d",
          9198 => x"69",
          9199 => x"05",
          9200 => x"72",
          9201 => x"5c",
          9202 => x"59",
          9203 => x"2e",
          9204 => x"89",
          9205 => x"60",
          9206 => x"84",
          9207 => x"5d",
          9208 => x"18",
          9209 => x"68",
          9210 => x"74",
          9211 => x"af",
          9212 => x"31",
          9213 => x"53",
          9214 => x"52",
          9215 => x"b1",
          9216 => x"d8",
          9217 => x"83",
          9218 => x"06",
          9219 => x"d6",
          9220 => x"ff",
          9221 => x"dd",
          9222 => x"83",
          9223 => x"2a",
          9224 => x"be",
          9225 => x"39",
          9226 => x"09",
          9227 => x"c5",
          9228 => x"f5",
          9229 => x"d8",
          9230 => x"38",
          9231 => x"79",
          9232 => x"80",
          9233 => x"38",
          9234 => x"96",
          9235 => x"06",
          9236 => x"2e",
          9237 => x"5e",
          9238 => x"82",
          9239 => x"9f",
          9240 => x"38",
          9241 => x"38",
          9242 => x"81",
          9243 => x"fc",
          9244 => x"ab",
          9245 => x"7d",
          9246 => x"81",
          9247 => x"7d",
          9248 => x"78",
          9249 => x"74",
          9250 => x"8e",
          9251 => x"9c",
          9252 => x"53",
          9253 => x"51",
          9254 => x"3f",
          9255 => x"c7",
          9256 => x"51",
          9257 => x"3f",
          9258 => x"8b",
          9259 => x"8f",
          9260 => x"8d",
          9261 => x"83",
          9262 => x"52",
          9263 => x"ff",
          9264 => x"81",
          9265 => x"34",
          9266 => x"70",
          9267 => x"2a",
          9268 => x"54",
          9269 => x"1b",
          9270 => x"b6",
          9271 => x"74",
          9272 => x"26",
          9273 => x"83",
          9274 => x"52",
          9275 => x"ff",
          9276 => x"8a",
          9277 => x"a0",
          9278 => x"8f",
          9279 => x"0b",
          9280 => x"bf",
          9281 => x"51",
          9282 => x"3f",
          9283 => x"9a",
          9284 => x"8e",
          9285 => x"52",
          9286 => x"ff",
          9287 => x"7d",
          9288 => x"81",
          9289 => x"38",
          9290 => x"0a",
          9291 => x"1b",
          9292 => x"fc",
          9293 => x"a4",
          9294 => x"8e",
          9295 => x"52",
          9296 => x"ff",
          9297 => x"81",
          9298 => x"51",
          9299 => x"3f",
          9300 => x"1b",
          9301 => x"ba",
          9302 => x"0b",
          9303 => x"34",
          9304 => x"c2",
          9305 => x"53",
          9306 => x"52",
          9307 => x"51",
          9308 => x"88",
          9309 => x"a7",
          9310 => x"8e",
          9311 => x"83",
          9312 => x"52",
          9313 => x"ff",
          9314 => x"ff",
          9315 => x"1c",
          9316 => x"a6",
          9317 => x"53",
          9318 => x"52",
          9319 => x"ff",
          9320 => x"82",
          9321 => x"83",
          9322 => x"52",
          9323 => x"e2",
          9324 => x"60",
          9325 => x"7e",
          9326 => x"85",
          9327 => x"82",
          9328 => x"83",
          9329 => x"83",
          9330 => x"06",
          9331 => x"75",
          9332 => x"05",
          9333 => x"7e",
          9334 => x"e5",
          9335 => x"53",
          9336 => x"51",
          9337 => x"3f",
          9338 => x"a4",
          9339 => x"51",
          9340 => x"3f",
          9341 => x"e4",
          9342 => x"e4",
          9343 => x"8d",
          9344 => x"18",
          9345 => x"1b",
          9346 => x"a4",
          9347 => x"83",
          9348 => x"ff",
          9349 => x"82",
          9350 => x"78",
          9351 => x"f2",
          9352 => x"60",
          9353 => x"7a",
          9354 => x"ff",
          9355 => x"75",
          9356 => x"53",
          9357 => x"51",
          9358 => x"3f",
          9359 => x"52",
          9360 => x"8d",
          9361 => x"56",
          9362 => x"83",
          9363 => x"06",
          9364 => x"52",
          9365 => x"8c",
          9366 => x"52",
          9367 => x"ff",
          9368 => x"f0",
          9369 => x"1b",
          9370 => x"87",
          9371 => x"55",
          9372 => x"83",
          9373 => x"74",
          9374 => x"ff",
          9375 => x"7c",
          9376 => x"74",
          9377 => x"38",
          9378 => x"54",
          9379 => x"52",
          9380 => x"88",
          9381 => x"d6",
          9382 => x"87",
          9383 => x"53",
          9384 => x"08",
          9385 => x"ff",
          9386 => x"76",
          9387 => x"31",
          9388 => x"cd",
          9389 => x"58",
          9390 => x"ff",
          9391 => x"55",
          9392 => x"83",
          9393 => x"61",
          9394 => x"26",
          9395 => x"57",
          9396 => x"53",
          9397 => x"51",
          9398 => x"3f",
          9399 => x"08",
          9400 => x"76",
          9401 => x"31",
          9402 => x"db",
          9403 => x"7d",
          9404 => x"38",
          9405 => x"83",
          9406 => x"8a",
          9407 => x"7d",
          9408 => x"38",
          9409 => x"81",
          9410 => x"80",
          9411 => x"80",
          9412 => x"7a",
          9413 => x"ea",
          9414 => x"d5",
          9415 => x"ff",
          9416 => x"83",
          9417 => x"77",
          9418 => x"0b",
          9419 => x"81",
          9420 => x"34",
          9421 => x"34",
          9422 => x"34",
          9423 => x"56",
          9424 => x"52",
          9425 => x"a1",
          9426 => x"0b",
          9427 => x"82",
          9428 => x"82",
          9429 => x"56",
          9430 => x"34",
          9431 => x"08",
          9432 => x"60",
          9433 => x"1b",
          9434 => x"c4",
          9435 => x"83",
          9436 => x"ff",
          9437 => x"81",
          9438 => x"7a",
          9439 => x"ff",
          9440 => x"81",
          9441 => x"d8",
          9442 => x"80",
          9443 => x"7e",
          9444 => x"91",
          9445 => x"82",
          9446 => x"90",
          9447 => x"8e",
          9448 => x"81",
          9449 => x"82",
          9450 => x"56",
          9451 => x"d8",
          9452 => x"0d",
          9453 => x"0d",
          9454 => x"59",
          9455 => x"ff",
          9456 => x"57",
          9457 => x"b4",
          9458 => x"f8",
          9459 => x"81",
          9460 => x"52",
          9461 => x"bd",
          9462 => x"2e",
          9463 => x"9c",
          9464 => x"33",
          9465 => x"2e",
          9466 => x"76",
          9467 => x"58",
          9468 => x"57",
          9469 => x"09",
          9470 => x"38",
          9471 => x"78",
          9472 => x"38",
          9473 => x"82",
          9474 => x"8d",
          9475 => x"f7",
          9476 => x"02",
          9477 => x"05",
          9478 => x"77",
          9479 => x"81",
          9480 => x"8d",
          9481 => x"e7",
          9482 => x"08",
          9483 => x"24",
          9484 => x"17",
          9485 => x"8c",
          9486 => x"77",
          9487 => x"16",
          9488 => x"25",
          9489 => x"3d",
          9490 => x"75",
          9491 => x"52",
          9492 => x"cb",
          9493 => x"76",
          9494 => x"70",
          9495 => x"2a",
          9496 => x"51",
          9497 => x"84",
          9498 => x"19",
          9499 => x"8b",
          9500 => x"f9",
          9501 => x"84",
          9502 => x"56",
          9503 => x"a7",
          9504 => x"fc",
          9505 => x"53",
          9506 => x"75",
          9507 => x"85",
          9508 => x"d8",
          9509 => x"84",
          9510 => x"2e",
          9511 => x"87",
          9512 => x"08",
          9513 => x"ff",
          9514 => x"d6",
          9515 => x"3d",
          9516 => x"3d",
          9517 => x"80",
          9518 => x"52",
          9519 => x"88",
          9520 => x"74",
          9521 => x"0d",
          9522 => x"0d",
          9523 => x"05",
          9524 => x"86",
          9525 => x"54",
          9526 => x"73",
          9527 => x"fe",
          9528 => x"51",
          9529 => x"98",
          9530 => x"fd",
          9531 => x"02",
          9532 => x"05",
          9533 => x"80",
          9534 => x"ff",
          9535 => x"72",
          9536 => x"06",
          9537 => x"39",
          9538 => x"73",
          9539 => x"83",
          9540 => x"81",
          9541 => x"70",
          9542 => x"38",
          9543 => x"22",
          9544 => x"2e",
          9545 => x"12",
          9546 => x"ff",
          9547 => x"71",
          9548 => x"8d",
          9549 => x"82",
          9550 => x"70",
          9551 => x"e1",
          9552 => x"12",
          9553 => x"06",
          9554 => x"82",
          9555 => x"85",
          9556 => x"fe",
          9557 => x"92",
          9558 => x"84",
          9559 => x"22",
          9560 => x"53",
          9561 => x"26",
          9562 => x"53",
          9563 => x"83",
          9564 => x"81",
          9565 => x"70",
          9566 => x"8b",
          9567 => x"82",
          9568 => x"70",
          9569 => x"72",
          9570 => x"0c",
          9571 => x"04",
          9572 => x"77",
          9573 => x"ff",
          9574 => x"a7",
          9575 => x"ff",
          9576 => x"cb",
          9577 => x"9f",
          9578 => x"85",
          9579 => x"8c",
          9580 => x"82",
          9581 => x"70",
          9582 => x"25",
          9583 => x"07",
          9584 => x"70",
          9585 => x"75",
          9586 => x"57",
          9587 => x"2a",
          9588 => x"06",
          9589 => x"52",
          9590 => x"71",
          9591 => x"38",
          9592 => x"80",
          9593 => x"84",
          9594 => x"98",
          9595 => x"08",
          9596 => x"31",
          9597 => x"70",
          9598 => x"51",
          9599 => x"71",
          9600 => x"06",
          9601 => x"51",
          9602 => x"f0",
          9603 => x"39",
          9604 => x"9a",
          9605 => x"51",
          9606 => x"12",
          9607 => x"88",
          9608 => x"39",
          9609 => x"51",
          9610 => x"a0",
          9611 => x"83",
          9612 => x"52",
          9613 => x"fe",
          9614 => x"10",
          9615 => x"f1",
          9616 => x"70",
          9617 => x"0c",
          9618 => x"04",
          9619 => x"00",
          9620 => x"ff",
          9621 => x"ff",
          9622 => x"ff",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"64",
          9769 => x"74",
          9770 => x"64",
          9771 => x"74",
          9772 => x"66",
          9773 => x"74",
          9774 => x"66",
          9775 => x"64",
          9776 => x"66",
          9777 => x"63",
          9778 => x"6d",
          9779 => x"61",
          9780 => x"6d",
          9781 => x"79",
          9782 => x"6d",
          9783 => x"66",
          9784 => x"6d",
          9785 => x"70",
          9786 => x"6d",
          9787 => x"6d",
          9788 => x"6d",
          9789 => x"68",
          9790 => x"68",
          9791 => x"68",
          9792 => x"68",
          9793 => x"63",
          9794 => x"00",
          9795 => x"6a",
          9796 => x"72",
          9797 => x"61",
          9798 => x"72",
          9799 => x"74",
          9800 => x"69",
          9801 => x"00",
          9802 => x"74",
          9803 => x"00",
          9804 => x"74",
          9805 => x"69",
          9806 => x"6d",
          9807 => x"69",
          9808 => x"6b",
          9809 => x"00",
          9810 => x"65",
          9811 => x"44",
          9812 => x"20",
          9813 => x"6f",
          9814 => x"49",
          9815 => x"72",
          9816 => x"20",
          9817 => x"6f",
          9818 => x"44",
          9819 => x"20",
          9820 => x"20",
          9821 => x"64",
          9822 => x"4e",
          9823 => x"69",
          9824 => x"66",
          9825 => x"64",
          9826 => x"4e",
          9827 => x"61",
          9828 => x"66",
          9829 => x"64",
          9830 => x"49",
          9831 => x"6c",
          9832 => x"66",
          9833 => x"6e",
          9834 => x"2e",
          9835 => x"41",
          9836 => x"73",
          9837 => x"65",
          9838 => x"64",
          9839 => x"46",
          9840 => x"20",
          9841 => x"65",
          9842 => x"20",
          9843 => x"73",
          9844 => x"00",
          9845 => x"46",
          9846 => x"20",
          9847 => x"64",
          9848 => x"69",
          9849 => x"6c",
          9850 => x"00",
          9851 => x"53",
          9852 => x"73",
          9853 => x"69",
          9854 => x"70",
          9855 => x"65",
          9856 => x"64",
          9857 => x"44",
          9858 => x"65",
          9859 => x"6d",
          9860 => x"20",
          9861 => x"69",
          9862 => x"6c",
          9863 => x"00",
          9864 => x"44",
          9865 => x"20",
          9866 => x"20",
          9867 => x"62",
          9868 => x"2e",
          9869 => x"4e",
          9870 => x"6f",
          9871 => x"74",
          9872 => x"65",
          9873 => x"6c",
          9874 => x"73",
          9875 => x"20",
          9876 => x"6e",
          9877 => x"6e",
          9878 => x"73",
          9879 => x"46",
          9880 => x"61",
          9881 => x"62",
          9882 => x"65",
          9883 => x"54",
          9884 => x"6f",
          9885 => x"20",
          9886 => x"72",
          9887 => x"6f",
          9888 => x"61",
          9889 => x"6c",
          9890 => x"2e",
          9891 => x"46",
          9892 => x"20",
          9893 => x"6c",
          9894 => x"65",
          9895 => x"49",
          9896 => x"66",
          9897 => x"69",
          9898 => x"20",
          9899 => x"6f",
          9900 => x"00",
          9901 => x"54",
          9902 => x"6d",
          9903 => x"20",
          9904 => x"6e",
          9905 => x"6c",
          9906 => x"00",
          9907 => x"50",
          9908 => x"6d",
          9909 => x"72",
          9910 => x"6e",
          9911 => x"72",
          9912 => x"2e",
          9913 => x"53",
          9914 => x"65",
          9915 => x"00",
          9916 => x"55",
          9917 => x"6f",
          9918 => x"65",
          9919 => x"72",
          9920 => x"0a",
          9921 => x"20",
          9922 => x"65",
          9923 => x"73",
          9924 => x"20",
          9925 => x"20",
          9926 => x"65",
          9927 => x"65",
          9928 => x"00",
          9929 => x"72",
          9930 => x"00",
          9931 => x"30",
          9932 => x"38",
          9933 => x"20",
          9934 => x"30",
          9935 => x"2c",
          9936 => x"25",
          9937 => x"78",
          9938 => x"49",
          9939 => x"25",
          9940 => x"78",
          9941 => x"38",
          9942 => x"25",
          9943 => x"78",
          9944 => x"25",
          9945 => x"58",
          9946 => x"3a",
          9947 => x"25",
          9948 => x"00",
          9949 => x"20",
          9950 => x"20",
          9951 => x"00",
          9952 => x"25",
          9953 => x"00",
          9954 => x"20",
          9955 => x"20",
          9956 => x"7c",
          9957 => x"7a",
          9958 => x"0a",
          9959 => x"25",
          9960 => x"00",
          9961 => x"30",
          9962 => x"32",
          9963 => x"32",
          9964 => x"76",
          9965 => x"34",
          9966 => x"20",
          9967 => x"2c",
          9968 => x"76",
          9969 => x"32",
          9970 => x"25",
          9971 => x"73",
          9972 => x"0a",
          9973 => x"5a",
          9974 => x"49",
          9975 => x"72",
          9976 => x"74",
          9977 => x"6e",
          9978 => x"72",
          9979 => x"54",
          9980 => x"72",
          9981 => x"74",
          9982 => x"75",
          9983 => x"50",
          9984 => x"69",
          9985 => x"72",
          9986 => x"74",
          9987 => x"49",
          9988 => x"4c",
          9989 => x"20",
          9990 => x"65",
          9991 => x"70",
          9992 => x"49",
          9993 => x"4c",
          9994 => x"20",
          9995 => x"65",
          9996 => x"70",
          9997 => x"55",
          9998 => x"30",
          9999 => x"20",
         10000 => x"65",
         10001 => x"70",
         10002 => x"55",
         10003 => x"30",
         10004 => x"20",
         10005 => x"65",
         10006 => x"70",
         10007 => x"55",
         10008 => x"31",
         10009 => x"20",
         10010 => x"65",
         10011 => x"70",
         10012 => x"55",
         10013 => x"31",
         10014 => x"20",
         10015 => x"65",
         10016 => x"70",
         10017 => x"53",
         10018 => x"69",
         10019 => x"75",
         10020 => x"69",
         10021 => x"2e",
         10022 => x"45",
         10023 => x"6c",
         10024 => x"20",
         10025 => x"65",
         10026 => x"2e",
         10027 => x"61",
         10028 => x"65",
         10029 => x"2e",
         10030 => x"00",
         10031 => x"7a",
         10032 => x"68",
         10033 => x"30",
         10034 => x"46",
         10035 => x"65",
         10036 => x"6f",
         10037 => x"69",
         10038 => x"6c",
         10039 => x"20",
         10040 => x"63",
         10041 => x"20",
         10042 => x"70",
         10043 => x"73",
         10044 => x"6e",
         10045 => x"6d",
         10046 => x"61",
         10047 => x"2e",
         10048 => x"2a",
         10049 => x"43",
         10050 => x"72",
         10051 => x"2e",
         10052 => x"00",
         10053 => x"43",
         10054 => x"69",
         10055 => x"2e",
         10056 => x"43",
         10057 => x"61",
         10058 => x"67",
         10059 => x"00",
         10060 => x"25",
         10061 => x"78",
         10062 => x"38",
         10063 => x"3e",
         10064 => x"6c",
         10065 => x"30",
         10066 => x"0a",
         10067 => x"44",
         10068 => x"20",
         10069 => x"6f",
         10070 => x"0a",
         10071 => x"70",
         10072 => x"65",
         10073 => x"25",
         10074 => x"58",
         10075 => x"32",
         10076 => x"3f",
         10077 => x"25",
         10078 => x"58",
         10079 => x"34",
         10080 => x"25",
         10081 => x"58",
         10082 => x"38",
         10083 => x"00",
         10084 => x"45",
         10085 => x"75",
         10086 => x"67",
         10087 => x"64",
         10088 => x"20",
         10089 => x"6c",
         10090 => x"2e",
         10091 => x"43",
         10092 => x"69",
         10093 => x"63",
         10094 => x"20",
         10095 => x"30",
         10096 => x"20",
         10097 => x"0a",
         10098 => x"43",
         10099 => x"20",
         10100 => x"75",
         10101 => x"64",
         10102 => x"64",
         10103 => x"25",
         10104 => x"0a",
         10105 => x"52",
         10106 => x"61",
         10107 => x"6e",
         10108 => x"70",
         10109 => x"63",
         10110 => x"6f",
         10111 => x"2e",
         10112 => x"43",
         10113 => x"20",
         10114 => x"6f",
         10115 => x"6e",
         10116 => x"2e",
         10117 => x"5a",
         10118 => x"62",
         10119 => x"25",
         10120 => x"25",
         10121 => x"73",
         10122 => x"00",
         10123 => x"25",
         10124 => x"25",
         10125 => x"73",
         10126 => x"25",
         10127 => x"25",
         10128 => x"42",
         10129 => x"63",
         10130 => x"61",
         10131 => x"00",
         10132 => x"4d",
         10133 => x"72",
         10134 => x"78",
         10135 => x"73",
         10136 => x"2c",
         10137 => x"6e",
         10138 => x"20",
         10139 => x"63",
         10140 => x"20",
         10141 => x"6d",
         10142 => x"2e",
         10143 => x"54",
         10144 => x"69",
         10145 => x"70",
         10146 => x"74",
         10147 => x"52",
         10148 => x"69",
         10149 => x"2e",
         10150 => x"45",
         10151 => x"6c",
         10152 => x"20",
         10153 => x"65",
         10154 => x"70",
         10155 => x"2e",
         10156 => x"25",
         10157 => x"64",
         10158 => x"20",
         10159 => x"25",
         10160 => x"64",
         10161 => x"25",
         10162 => x"53",
         10163 => x"43",
         10164 => x"69",
         10165 => x"61",
         10166 => x"6e",
         10167 => x"20",
         10168 => x"6f",
         10169 => x"6f",
         10170 => x"6f",
         10171 => x"67",
         10172 => x"3a",
         10173 => x"76",
         10174 => x"73",
         10175 => x"70",
         10176 => x"65",
         10177 => x"64",
         10178 => x"20",
         10179 => x"57",
         10180 => x"44",
         10181 => x"20",
         10182 => x"30",
         10183 => x"25",
         10184 => x"29",
         10185 => x"20",
         10186 => x"53",
         10187 => x"4d",
         10188 => x"20",
         10189 => x"30",
         10190 => x"25",
         10191 => x"29",
         10192 => x"20",
         10193 => x"49",
         10194 => x"20",
         10195 => x"4d",
         10196 => x"30",
         10197 => x"25",
         10198 => x"29",
         10199 => x"20",
         10200 => x"42",
         10201 => x"20",
         10202 => x"20",
         10203 => x"30",
         10204 => x"25",
         10205 => x"29",
         10206 => x"20",
         10207 => x"52",
         10208 => x"20",
         10209 => x"20",
         10210 => x"30",
         10211 => x"25",
         10212 => x"29",
         10213 => x"20",
         10214 => x"53",
         10215 => x"41",
         10216 => x"20",
         10217 => x"65",
         10218 => x"65",
         10219 => x"25",
         10220 => x"29",
         10221 => x"20",
         10222 => x"54",
         10223 => x"52",
         10224 => x"20",
         10225 => x"69",
         10226 => x"73",
         10227 => x"25",
         10228 => x"29",
         10229 => x"20",
         10230 => x"49",
         10231 => x"20",
         10232 => x"4c",
         10233 => x"68",
         10234 => x"65",
         10235 => x"25",
         10236 => x"29",
         10237 => x"20",
         10238 => x"57",
         10239 => x"42",
         10240 => x"20",
         10241 => x"00",
         10242 => x"20",
         10243 => x"57",
         10244 => x"32",
         10245 => x"20",
         10246 => x"49",
         10247 => x"4c",
         10248 => x"20",
         10249 => x"50",
         10250 => x"20",
         10251 => x"53",
         10252 => x"41",
         10253 => x"65",
         10254 => x"73",
         10255 => x"20",
         10256 => x"43",
         10257 => x"52",
         10258 => x"74",
         10259 => x"63",
         10260 => x"20",
         10261 => x"72",
         10262 => x"20",
         10263 => x"30",
         10264 => x"00",
         10265 => x"20",
         10266 => x"43",
         10267 => x"4d",
         10268 => x"72",
         10269 => x"74",
         10270 => x"20",
         10271 => x"72",
         10272 => x"20",
         10273 => x"30",
         10274 => x"00",
         10275 => x"20",
         10276 => x"53",
         10277 => x"6b",
         10278 => x"61",
         10279 => x"41",
         10280 => x"65",
         10281 => x"20",
         10282 => x"20",
         10283 => x"30",
         10284 => x"00",
         10285 => x"4d",
         10286 => x"3a",
         10287 => x"20",
         10288 => x"5a",
         10289 => x"49",
         10290 => x"20",
         10291 => x"20",
         10292 => x"20",
         10293 => x"20",
         10294 => x"20",
         10295 => x"30",
         10296 => x"00",
         10297 => x"20",
         10298 => x"53",
         10299 => x"65",
         10300 => x"6c",
         10301 => x"20",
         10302 => x"71",
         10303 => x"20",
         10304 => x"20",
         10305 => x"64",
         10306 => x"34",
         10307 => x"7a",
         10308 => x"20",
         10309 => x"53",
         10310 => x"4d",
         10311 => x"6f",
         10312 => x"46",
         10313 => x"20",
         10314 => x"20",
         10315 => x"20",
         10316 => x"64",
         10317 => x"34",
         10318 => x"7a",
         10319 => x"20",
         10320 => x"57",
         10321 => x"62",
         10322 => x"20",
         10323 => x"41",
         10324 => x"6c",
         10325 => x"20",
         10326 => x"71",
         10327 => x"64",
         10328 => x"34",
         10329 => x"7a",
         10330 => x"53",
         10331 => x"6c",
         10332 => x"4d",
         10333 => x"75",
         10334 => x"46",
         10335 => x"00",
         10336 => x"45",
         10337 => x"45",
         10338 => x"00",
         10339 => x"55",
         10340 => x"6f",
         10341 => x"00",
         10342 => x"01",
         10343 => x"00",
         10344 => x"00",
         10345 => x"01",
         10346 => x"00",
         10347 => x"00",
         10348 => x"01",
         10349 => x"00",
         10350 => x"00",
         10351 => x"01",
         10352 => x"00",
         10353 => x"00",
         10354 => x"01",
         10355 => x"00",
         10356 => x"00",
         10357 => x"01",
         10358 => x"00",
         10359 => x"00",
         10360 => x"01",
         10361 => x"00",
         10362 => x"00",
         10363 => x"01",
         10364 => x"00",
         10365 => x"00",
         10366 => x"01",
         10367 => x"00",
         10368 => x"00",
         10369 => x"01",
         10370 => x"00",
         10371 => x"00",
         10372 => x"01",
         10373 => x"00",
         10374 => x"00",
         10375 => x"04",
         10376 => x"00",
         10377 => x"00",
         10378 => x"04",
         10379 => x"00",
         10380 => x"00",
         10381 => x"04",
         10382 => x"00",
         10383 => x"00",
         10384 => x"03",
         10385 => x"00",
         10386 => x"00",
         10387 => x"04",
         10388 => x"00",
         10389 => x"00",
         10390 => x"04",
         10391 => x"00",
         10392 => x"00",
         10393 => x"04",
         10394 => x"00",
         10395 => x"00",
         10396 => x"03",
         10397 => x"00",
         10398 => x"00",
         10399 => x"03",
         10400 => x"00",
         10401 => x"00",
         10402 => x"03",
         10403 => x"00",
         10404 => x"00",
         10405 => x"03",
         10406 => x"00",
         10407 => x"1b",
         10408 => x"1b",
         10409 => x"1b",
         10410 => x"1b",
         10411 => x"1b",
         10412 => x"1b",
         10413 => x"1b",
         10414 => x"1b",
         10415 => x"1b",
         10416 => x"1b",
         10417 => x"1b",
         10418 => x"10",
         10419 => x"0e",
         10420 => x"0d",
         10421 => x"0b",
         10422 => x"08",
         10423 => x"06",
         10424 => x"05",
         10425 => x"04",
         10426 => x"03",
         10427 => x"02",
         10428 => x"01",
         10429 => x"68",
         10430 => x"6f",
         10431 => x"68",
         10432 => x"00",
         10433 => x"21",
         10434 => x"25",
         10435 => x"75",
         10436 => x"73",
         10437 => x"46",
         10438 => x"65",
         10439 => x"6f",
         10440 => x"73",
         10441 => x"74",
         10442 => x"68",
         10443 => x"6f",
         10444 => x"66",
         10445 => x"20",
         10446 => x"45",
         10447 => x"00",
         10448 => x"43",
         10449 => x"6f",
         10450 => x"70",
         10451 => x"63",
         10452 => x"74",
         10453 => x"69",
         10454 => x"72",
         10455 => x"69",
         10456 => x"20",
         10457 => x"61",
         10458 => x"6e",
         10459 => x"53",
         10460 => x"22",
         10461 => x"3e",
         10462 => x"00",
         10463 => x"2b",
         10464 => x"5b",
         10465 => x"46",
         10466 => x"46",
         10467 => x"32",
         10468 => x"eb",
         10469 => x"53",
         10470 => x"35",
         10471 => x"4e",
         10472 => x"41",
         10473 => x"20",
         10474 => x"41",
         10475 => x"20",
         10476 => x"4e",
         10477 => x"41",
         10478 => x"20",
         10479 => x"41",
         10480 => x"20",
         10481 => x"00",
         10482 => x"00",
         10483 => x"00",
         10484 => x"00",
         10485 => x"01",
         10486 => x"09",
         10487 => x"14",
         10488 => x"1e",
         10489 => x"80",
         10490 => x"8e",
         10491 => x"45",
         10492 => x"49",
         10493 => x"90",
         10494 => x"99",
         10495 => x"59",
         10496 => x"9c",
         10497 => x"41",
         10498 => x"a5",
         10499 => x"a8",
         10500 => x"ac",
         10501 => x"b0",
         10502 => x"b4",
         10503 => x"b8",
         10504 => x"bc",
         10505 => x"c0",
         10506 => x"c4",
         10507 => x"c8",
         10508 => x"cc",
         10509 => x"d0",
         10510 => x"d4",
         10511 => x"d8",
         10512 => x"dc",
         10513 => x"e0",
         10514 => x"e4",
         10515 => x"e8",
         10516 => x"ec",
         10517 => x"f0",
         10518 => x"f4",
         10519 => x"f8",
         10520 => x"fc",
         10521 => x"2b",
         10522 => x"3d",
         10523 => x"5c",
         10524 => x"3c",
         10525 => x"7f",
         10526 => x"00",
         10527 => x"00",
         10528 => x"01",
         10529 => x"00",
         10530 => x"00",
         10531 => x"00",
         10532 => x"00",
         10533 => x"00",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"00",
         10538 => x"00",
         10539 => x"00",
         10540 => x"00",
         10541 => x"00",
         10542 => x"00",
         10543 => x"00",
         10544 => x"00",
         10545 => x"00",
         10546 => x"00",
         10547 => x"00",
         10548 => x"00",
         10549 => x"20",
         10550 => x"00",
         10551 => x"00",
         10552 => x"00",
         10553 => x"00",
         10554 => x"00",
         10555 => x"00",
         10556 => x"00",
         10557 => x"00",
         10558 => x"25",
         10559 => x"25",
         10560 => x"25",
         10561 => x"25",
         10562 => x"25",
         10563 => x"25",
         10564 => x"25",
         10565 => x"25",
         10566 => x"25",
         10567 => x"25",
         10568 => x"25",
         10569 => x"25",
         10570 => x"25",
         10571 => x"25",
         10572 => x"25",
         10573 => x"25",
         10574 => x"25",
         10575 => x"25",
         10576 => x"25",
         10577 => x"25",
         10578 => x"25",
         10579 => x"25",
         10580 => x"25",
         10581 => x"25",
         10582 => x"03",
         10583 => x"03",
         10584 => x"03",
         10585 => x"00",
         10586 => x"03",
         10587 => x"03",
         10588 => x"22",
         10589 => x"03",
         10590 => x"22",
         10591 => x"22",
         10592 => x"23",
         10593 => x"00",
         10594 => x"00",
         10595 => x"00",
         10596 => x"20",
         10597 => x"25",
         10598 => x"00",
         10599 => x"00",
         10600 => x"00",
         10601 => x"00",
         10602 => x"01",
         10603 => x"01",
         10604 => x"01",
         10605 => x"01",
         10606 => x"01",
         10607 => x"01",
         10608 => x"00",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"01",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"01",
         10622 => x"01",
         10623 => x"01",
         10624 => x"01",
         10625 => x"01",
         10626 => x"01",
         10627 => x"01",
         10628 => x"01",
         10629 => x"01",
         10630 => x"01",
         10631 => x"01",
         10632 => x"01",
         10633 => x"01",
         10634 => x"01",
         10635 => x"01",
         10636 => x"01",
         10637 => x"01",
         10638 => x"01",
         10639 => x"01",
         10640 => x"01",
         10641 => x"01",
         10642 => x"01",
         10643 => x"01",
         10644 => x"01",
         10645 => x"01",
         10646 => x"01",
         10647 => x"01",
         10648 => x"01",
         10649 => x"01",
         10650 => x"01",
         10651 => x"00",
         10652 => x"01",
         10653 => x"01",
         10654 => x"02",
         10655 => x"02",
         10656 => x"2c",
         10657 => x"02",
         10658 => x"2c",
         10659 => x"02",
         10660 => x"02",
         10661 => x"01",
         10662 => x"00",
         10663 => x"01",
         10664 => x"01",
         10665 => x"02",
         10666 => x"02",
         10667 => x"02",
         10668 => x"02",
         10669 => x"01",
         10670 => x"02",
         10671 => x"02",
         10672 => x"02",
         10673 => x"01",
         10674 => x"02",
         10675 => x"02",
         10676 => x"02",
         10677 => x"02",
         10678 => x"01",
         10679 => x"02",
         10680 => x"02",
         10681 => x"02",
         10682 => x"02",
         10683 => x"02",
         10684 => x"02",
         10685 => x"01",
         10686 => x"02",
         10687 => x"02",
         10688 => x"02",
         10689 => x"01",
         10690 => x"01",
         10691 => x"02",
         10692 => x"02",
         10693 => x"02",
         10694 => x"01",
         10695 => x"00",
         10696 => x"03",
         10697 => x"03",
         10698 => x"03",
         10699 => x"03",
         10700 => x"03",
         10701 => x"03",
         10702 => x"03",
         10703 => x"03",
         10704 => x"03",
         10705 => x"03",
         10706 => x"03",
         10707 => x"01",
         10708 => x"00",
         10709 => x"03",
         10710 => x"03",
         10711 => x"03",
         10712 => x"03",
         10713 => x"03",
         10714 => x"03",
         10715 => x"07",
         10716 => x"01",
         10717 => x"01",
         10718 => x"01",
         10719 => x"00",
         10720 => x"04",
         10721 => x"05",
         10722 => x"00",
         10723 => x"1d",
         10724 => x"2c",
         10725 => x"01",
         10726 => x"01",
         10727 => x"06",
         10728 => x"06",
         10729 => x"06",
         10730 => x"06",
         10731 => x"06",
         10732 => x"00",
         10733 => x"1f",
         10734 => x"1f",
         10735 => x"1f",
         10736 => x"1f",
         10737 => x"1f",
         10738 => x"1f",
         10739 => x"1f",
         10740 => x"1f",
         10741 => x"1f",
         10742 => x"1f",
         10743 => x"1f",
         10744 => x"1f",
         10745 => x"1f",
         10746 => x"1f",
         10747 => x"1f",
         10748 => x"1f",
         10749 => x"1f",
         10750 => x"1f",
         10751 => x"1f",
         10752 => x"1f",
         10753 => x"06",
         10754 => x"06",
         10755 => x"00",
         10756 => x"1f",
         10757 => x"1f",
         10758 => x"00",
         10759 => x"21",
         10760 => x"21",
         10761 => x"21",
         10762 => x"05",
         10763 => x"04",
         10764 => x"01",
         10765 => x"01",
         10766 => x"01",
         10767 => x"01",
         10768 => x"08",
         10769 => x"03",
         10770 => x"00",
         10771 => x"00",
         10772 => x"01",
         10773 => x"00",
         10774 => x"00",
         10775 => x"00",
         10776 => x"01",
         10777 => x"00",
         10778 => x"00",
         10779 => x"00",
         10780 => x"01",
         10781 => x"00",
         10782 => x"00",
         10783 => x"00",
         10784 => x"01",
         10785 => x"00",
         10786 => x"00",
         10787 => x"00",
         10788 => x"01",
         10789 => x"00",
         10790 => x"00",
         10791 => x"00",
         10792 => x"01",
         10793 => x"00",
         10794 => x"00",
         10795 => x"00",
         10796 => x"01",
         10797 => x"00",
         10798 => x"00",
         10799 => x"00",
         10800 => x"01",
         10801 => x"00",
         10802 => x"00",
         10803 => x"00",
         10804 => x"01",
         10805 => x"00",
         10806 => x"00",
         10807 => x"00",
         10808 => x"01",
         10809 => x"00",
         10810 => x"00",
         10811 => x"00",
         10812 => x"01",
         10813 => x"00",
         10814 => x"00",
         10815 => x"00",
         10816 => x"01",
         10817 => x"00",
         10818 => x"00",
         10819 => x"00",
         10820 => x"01",
         10821 => x"00",
         10822 => x"00",
         10823 => x"00",
         10824 => x"01",
         10825 => x"00",
         10826 => x"00",
         10827 => x"00",
         10828 => x"01",
         10829 => x"00",
         10830 => x"00",
         10831 => x"00",
         10832 => x"01",
         10833 => x"00",
         10834 => x"00",
         10835 => x"00",
         10836 => x"01",
         10837 => x"00",
         10838 => x"00",
         10839 => x"00",
         10840 => x"01",
         10841 => x"00",
         10842 => x"00",
         10843 => x"00",
         10844 => x"01",
         10845 => x"00",
         10846 => x"00",
         10847 => x"00",
         10848 => x"01",
         10849 => x"00",
         10850 => x"00",
         10851 => x"00",
         10852 => x"01",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"01",
         10857 => x"00",
         10858 => x"00",
         10859 => x"00",
         10860 => x"01",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"01",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"01",
         10869 => x"00",
         10870 => x"00",
         10871 => x"00",
         10872 => x"01",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"01",
         10885 => x"01",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"05",
         10891 => x"05",
         10892 => x"05",
         10893 => x"00",
         10894 => x"01",
         10895 => x"01",
         10896 => x"01",
         10897 => x"01",
         10898 => x"00",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"01",
         10924 => x"00",
         10925 => x"01",
         10926 => x"00",
         10927 => x"02",
         10928 => x"cc",
         10929 => x"ce",
         10930 => x"f8",
         10931 => x"fc",
         10932 => x"e1",
         10933 => x"c4",
         10934 => x"e3",
         10935 => x"eb",
         10936 => x"00",
         10937 => x"64",
         10938 => x"68",
         10939 => x"2f",
         10940 => x"20",
         10941 => x"24",
         10942 => x"28",
         10943 => x"51",
         10944 => x"55",
         10945 => x"04",
         10946 => x"08",
         10947 => x"0c",
         10948 => x"10",
         10949 => x"14",
         10950 => x"18",
         10951 => x"59",
         10952 => x"c7",
         10953 => x"84",
         10954 => x"88",
         10955 => x"8c",
         10956 => x"90",
         10957 => x"94",
         10958 => x"98",
         10959 => x"80",
         10960 => x"00",
         10961 => x"00",
         10962 => x"00",
         10963 => x"00",
         10964 => x"00",
         10965 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
