../../../../../cpu/zpu_core_evo_L2.vhd