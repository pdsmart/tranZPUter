-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b0b96",
          2049 => x"da040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b96",
          2121 => x"be040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b96a1",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81c4",
          2210 => x"d8738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"96a60400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b97",
          2219 => x"df2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b99",
          2227 => x"cb2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000800",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b90",
          2313 => x"81040b0b",
          2314 => x"0b908504",
          2315 => x"0b0b0b90",
          2316 => x"94040b0b",
          2317 => x"0b90a304",
          2318 => x"0b0b0b90",
          2319 => x"b2040b0b",
          2320 => x"0b90c104",
          2321 => x"0b0b0b90",
          2322 => x"d0040b0b",
          2323 => x"0b90df04",
          2324 => x"0b0b0b90",
          2325 => x"ee040b0b",
          2326 => x"0b90fd04",
          2327 => x"0b0b0b91",
          2328 => x"8c040b0b",
          2329 => x"0b919b04",
          2330 => x"0b0b0b91",
          2331 => x"aa040b0b",
          2332 => x"0b91b904",
          2333 => x"0b0b0b91",
          2334 => x"c8040b0b",
          2335 => x"0b91d704",
          2336 => x"0b0b0b91",
          2337 => x"e6040b0b",
          2338 => x"0b91f504",
          2339 => x"0b0b0b92",
          2340 => x"84040b0b",
          2341 => x"0b929404",
          2342 => x"0b0b0b92",
          2343 => x"a4040b0b",
          2344 => x"0b92b404",
          2345 => x"0b0b0b92",
          2346 => x"c4040b0b",
          2347 => x"0b92d404",
          2348 => x"0b0b0b92",
          2349 => x"e4040b0b",
          2350 => x"0b92f404",
          2351 => x"0b0b0b93",
          2352 => x"84040b0b",
          2353 => x"0b939404",
          2354 => x"0b0b0b93",
          2355 => x"a4040b0b",
          2356 => x"0b93b404",
          2357 => x"0b0b0b93",
          2358 => x"c4040b0b",
          2359 => x"0b93d404",
          2360 => x"0b0b0b93",
          2361 => x"e4040b0b",
          2362 => x"0b93f404",
          2363 => x"0b0b0b94",
          2364 => x"84040b0b",
          2365 => x"0b949404",
          2366 => x"0b0b0b94",
          2367 => x"a4040b0b",
          2368 => x"0b94b404",
          2369 => x"0b0b0b94",
          2370 => x"c4040b0b",
          2371 => x"0b94d404",
          2372 => x"0b0b0b94",
          2373 => x"e4040b0b",
          2374 => x"0b94f404",
          2375 => x"0b0b0b95",
          2376 => x"84040b0b",
          2377 => x"0b959404",
          2378 => x"0b0b0b95",
          2379 => x"a3040b0b",
          2380 => x"0b95b304",
          2381 => x"0b0b0b95",
          2382 => x"c3040b0b",
          2383 => x"0b95d204",
          2384 => x"0b0b0b95",
          2385 => x"e1040b0b",
          2386 => x"0b95f004",
          2387 => x"ffffffff",
          2388 => x"ffffffff",
          2389 => x"ffffffff",
          2390 => x"ffffffff",
          2391 => x"ffffffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"00000000",
          2433 => x"00000000",
          2434 => x"00000000",
          2435 => x"00000000",
          2436 => x"00000000",
          2437 => x"00000000",
          2438 => x"00000000",
          2439 => x"00000000",
          2440 => x"00000000",
          2441 => x"00000000",
          2442 => x"00000000",
          2443 => x"00000000",
          2444 => x"00000000",
          2445 => x"00000000",
          2446 => x"00000000",
          2447 => x"00000000",
          2448 => x"00000000",
          2449 => x"00000000",
          2450 => x"00000000",
          2451 => x"00000000",
          2452 => x"00000000",
          2453 => x"00000000",
          2454 => x"00000000",
          2455 => x"00000000",
          2456 => x"00000000",
          2457 => x"00000000",
          2458 => x"00000000",
          2459 => x"00000000",
          2460 => x"00000000",
          2461 => x"00000000",
          2462 => x"00000000",
          2463 => x"00000000",
          2464 => x"00000000",
          2465 => x"00000000",
          2466 => x"00000000",
          2467 => x"00000000",
          2468 => x"00000000",
          2469 => x"00000000",
          2470 => x"00000000",
          2471 => x"00000000",
          2472 => x"00000000",
          2473 => x"00000000",
          2474 => x"00000000",
          2475 => x"00000000",
          2476 => x"00000000",
          2477 => x"00000000",
          2478 => x"00000000",
          2479 => x"00000000",
          2480 => x"00000000",
          2481 => x"00000000",
          2482 => x"00000000",
          2483 => x"00000000",
          2484 => x"00000000",
          2485 => x"00000000",
          2486 => x"00000000",
          2487 => x"00000000",
          2488 => x"00000000",
          2489 => x"00000000",
          2490 => x"00000000",
          2491 => x"00000000",
          2492 => x"00000000",
          2493 => x"00000000",
          2494 => x"00000000",
          2495 => x"00000000",
          2496 => x"00000000",
          2497 => x"00000000",
          2498 => x"00000000",
          2499 => x"00000000",
          2500 => x"00000000",
          2501 => x"00000000",
          2502 => x"00000000",
          2503 => x"00000000",
          2504 => x"00000000",
          2505 => x"00000000",
          2506 => x"00000000",
          2507 => x"00000000",
          2508 => x"00000000",
          2509 => x"00000000",
          2510 => x"00000000",
          2511 => x"00000000",
          2512 => x"00000000",
          2513 => x"00000000",
          2514 => x"00000000",
          2515 => x"00000000",
          2516 => x"00000000",
          2517 => x"00000000",
          2518 => x"00000000",
          2519 => x"00000000",
          2520 => x"00000000",
          2521 => x"00000000",
          2522 => x"00000000",
          2523 => x"00000000",
          2524 => x"00000000",
          2525 => x"00000000",
          2526 => x"00000000",
          2527 => x"00000000",
          2528 => x"00000000",
          2529 => x"00000000",
          2530 => x"00000000",
          2531 => x"00000000",
          2532 => x"00000000",
          2533 => x"00000000",
          2534 => x"00000000",
          2535 => x"00000000",
          2536 => x"00000000",
          2537 => x"00000000",
          2538 => x"00000000",
          2539 => x"00000000",
          2540 => x"00000000",
          2541 => x"00000000",
          2542 => x"00000000",
          2543 => x"00000000",
          2544 => x"00000000",
          2545 => x"00000000",
          2546 => x"00000000",
          2547 => x"00000000",
          2548 => x"00000000",
          2549 => x"00000000",
          2550 => x"00000000",
          2551 => x"00000000",
          2552 => x"00000000",
          2553 => x"00000000",
          2554 => x"00000000",
          2555 => x"00000000",
          2556 => x"00000000",
          2557 => x"00000000",
          2558 => x"00000000",
          2559 => x"00000000",
          2560 => x"04009081",
          2561 => x"0481dcd8",
          2562 => x"0ca4b02d",
          2563 => x"81dcd808",
          2564 => x"83809004",
          2565 => x"81dcd80c",
          2566 => x"b1a32d81",
          2567 => x"dcd80883",
          2568 => x"80900481",
          2569 => x"dcd80cb1",
          2570 => x"e22d81dc",
          2571 => x"d8088380",
          2572 => x"900481dc",
          2573 => x"d80cb280",
          2574 => x"2d81dcd8",
          2575 => x"08838090",
          2576 => x"0481dcd8",
          2577 => x"0cb8be2d",
          2578 => x"81dcd808",
          2579 => x"83809004",
          2580 => x"81dcd80c",
          2581 => x"b9bc2d81",
          2582 => x"dcd80883",
          2583 => x"80900481",
          2584 => x"dcd80cb2",
          2585 => x"a32d81dc",
          2586 => x"d8088380",
          2587 => x"900481dc",
          2588 => x"d80cb9d9",
          2589 => x"2d81dcd8",
          2590 => x"08838090",
          2591 => x"0481dcd8",
          2592 => x"0cbbcb2d",
          2593 => x"81dcd808",
          2594 => x"83809004",
          2595 => x"81dcd80c",
          2596 => x"b7e42d81",
          2597 => x"dcd80883",
          2598 => x"80900481",
          2599 => x"dcd80cb7",
          2600 => x"fa2d81dc",
          2601 => x"d8088380",
          2602 => x"900481dc",
          2603 => x"d80cb89e",
          2604 => x"2d81dcd8",
          2605 => x"08838090",
          2606 => x"0481dcd8",
          2607 => x"0ca6bd2d",
          2608 => x"81dcd808",
          2609 => x"83809004",
          2610 => x"81dcd80c",
          2611 => x"a78e2d81",
          2612 => x"dcd80883",
          2613 => x"80900481",
          2614 => x"dcd80c9f",
          2615 => x"aa2d81dc",
          2616 => x"d8088380",
          2617 => x"900481dc",
          2618 => x"d80ca0df",
          2619 => x"2d81dcd8",
          2620 => x"08838090",
          2621 => x"0481dcd8",
          2622 => x"0ca2922d",
          2623 => x"81dcd808",
          2624 => x"83809004",
          2625 => x"81dcd80c",
          2626 => x"80ee802d",
          2627 => x"81dcd808",
          2628 => x"83809004",
          2629 => x"81dcd80c",
          2630 => x"80faf12d",
          2631 => x"81dcd808",
          2632 => x"83809004",
          2633 => x"81dcd80c",
          2634 => x"80f2e52d",
          2635 => x"81dcd808",
          2636 => x"83809004",
          2637 => x"81dcd80c",
          2638 => x"80f5e22d",
          2639 => x"81dcd808",
          2640 => x"83809004",
          2641 => x"81dcd80c",
          2642 => x"8180802d",
          2643 => x"81dcd808",
          2644 => x"83809004",
          2645 => x"81dcd80c",
          2646 => x"8188e02d",
          2647 => x"81dcd808",
          2648 => x"83809004",
          2649 => x"81dcd80c",
          2650 => x"80f9d32d",
          2651 => x"81dcd808",
          2652 => x"83809004",
          2653 => x"81dcd80c",
          2654 => x"81839f2d",
          2655 => x"81dcd808",
          2656 => x"83809004",
          2657 => x"81dcd80c",
          2658 => x"8184be2d",
          2659 => x"81dcd808",
          2660 => x"83809004",
          2661 => x"81dcd80c",
          2662 => x"8184dd2d",
          2663 => x"81dcd808",
          2664 => x"83809004",
          2665 => x"81dcd80c",
          2666 => x"818cc72d",
          2667 => x"81dcd808",
          2668 => x"83809004",
          2669 => x"81dcd80c",
          2670 => x"818aad2d",
          2671 => x"81dcd808",
          2672 => x"83809004",
          2673 => x"81dcd80c",
          2674 => x"818f9b2d",
          2675 => x"81dcd808",
          2676 => x"83809004",
          2677 => x"81dcd80c",
          2678 => x"8185e12d",
          2679 => x"81dcd808",
          2680 => x"83809004",
          2681 => x"81dcd80c",
          2682 => x"81929b2d",
          2683 => x"81dcd808",
          2684 => x"83809004",
          2685 => x"81dcd80c",
          2686 => x"81939c2d",
          2687 => x"81dcd808",
          2688 => x"83809004",
          2689 => x"81dcd80c",
          2690 => x"80fbd12d",
          2691 => x"81dcd808",
          2692 => x"83809004",
          2693 => x"81dcd80c",
          2694 => x"80fbaa2d",
          2695 => x"81dcd808",
          2696 => x"83809004",
          2697 => x"81dcd80c",
          2698 => x"80fcd52d",
          2699 => x"81dcd808",
          2700 => x"83809004",
          2701 => x"81dcd80c",
          2702 => x"8186b82d",
          2703 => x"81dcd808",
          2704 => x"83809004",
          2705 => x"81dcd80c",
          2706 => x"81948d2d",
          2707 => x"81dcd808",
          2708 => x"83809004",
          2709 => x"81dcd80c",
          2710 => x"8196972d",
          2711 => x"81dcd808",
          2712 => x"83809004",
          2713 => x"81dcd80c",
          2714 => x"8199d92d",
          2715 => x"81dcd808",
          2716 => x"83809004",
          2717 => x"81dcd80c",
          2718 => x"80ed9f2d",
          2719 => x"81dcd808",
          2720 => x"83809004",
          2721 => x"81dcd80c",
          2722 => x"819cc52d",
          2723 => x"81dcd808",
          2724 => x"83809004",
          2725 => x"81dcd80c",
          2726 => x"beda2d81",
          2727 => x"dcd80883",
          2728 => x"80900481",
          2729 => x"dcd80c80",
          2730 => x"c0c42d81",
          2731 => x"dcd80883",
          2732 => x"80900481",
          2733 => x"dcd80c80",
          2734 => x"c2a82d81",
          2735 => x"dcd80883",
          2736 => x"80900481",
          2737 => x"dcd80c9f",
          2738 => x"d32d81dc",
          2739 => x"d8088380",
          2740 => x"900481dc",
          2741 => x"d80ca0b5",
          2742 => x"2d81dcd8",
          2743 => x"08838090",
          2744 => x"0481dcd8",
          2745 => x"0ca3a22d",
          2746 => x"81dcd808",
          2747 => x"83809004",
          2748 => x"81dcd80c",
          2749 => x"81aac22d",
          2750 => x"81dcd808",
          2751 => x"83809004",
          2752 => x"3c041010",
          2753 => x"10101010",
          2754 => x"10101010",
          2755 => x"10101010",
          2756 => x"10101010",
          2757 => x"10101010",
          2758 => x"10101010",
          2759 => x"10101010",
          2760 => x"10535104",
          2761 => x"00007381",
          2762 => x"ff067383",
          2763 => x"06098105",
          2764 => x"83051010",
          2765 => x"102b0772",
          2766 => x"fc060c51",
          2767 => x"51047272",
          2768 => x"80728106",
          2769 => x"ff050972",
          2770 => x"06057110",
          2771 => x"52720a10",
          2772 => x"0a5372ed",
          2773 => x"38515153",
          2774 => x"510481dc",
          2775 => x"cc7081f3",
          2776 => x"f8278e38",
          2777 => x"80717084",
          2778 => x"05530c0b",
          2779 => x"0b0b96dd",
          2780 => x"04908151",
          2781 => x"81c3a704",
          2782 => x"0081dcd8",
          2783 => x"080281dc",
          2784 => x"d80cfd3d",
          2785 => x"0d805381",
          2786 => x"dcd8088c",
          2787 => x"05085281",
          2788 => x"dcd80888",
          2789 => x"05085183",
          2790 => x"d43f81dc",
          2791 => x"cc087081",
          2792 => x"dccc0c54",
          2793 => x"853d0d81",
          2794 => x"dcd80c04",
          2795 => x"81dcd808",
          2796 => x"0281dcd8",
          2797 => x"0cfd3d0d",
          2798 => x"815381dc",
          2799 => x"d8088c05",
          2800 => x"085281dc",
          2801 => x"d8088805",
          2802 => x"085183a1",
          2803 => x"3f81dccc",
          2804 => x"087081dc",
          2805 => x"cc0c5485",
          2806 => x"3d0d81dc",
          2807 => x"d80c0481",
          2808 => x"dcd80802",
          2809 => x"81dcd80c",
          2810 => x"f93d0d80",
          2811 => x"0b81dcd8",
          2812 => x"08fc050c",
          2813 => x"81dcd808",
          2814 => x"88050880",
          2815 => x"25b93881",
          2816 => x"dcd80888",
          2817 => x"05083081",
          2818 => x"dcd80888",
          2819 => x"050c800b",
          2820 => x"81dcd808",
          2821 => x"f4050c81",
          2822 => x"dcd808fc",
          2823 => x"05088a38",
          2824 => x"810b81dc",
          2825 => x"d808f405",
          2826 => x"0c81dcd8",
          2827 => x"08f40508",
          2828 => x"81dcd808",
          2829 => x"fc050c81",
          2830 => x"dcd8088c",
          2831 => x"05088025",
          2832 => x"b93881dc",
          2833 => x"d8088c05",
          2834 => x"083081dc",
          2835 => x"d8088c05",
          2836 => x"0c800b81",
          2837 => x"dcd808f0",
          2838 => x"050c81dc",
          2839 => x"d808fc05",
          2840 => x"088a3881",
          2841 => x"0b81dcd8",
          2842 => x"08f0050c",
          2843 => x"81dcd808",
          2844 => x"f0050881",
          2845 => x"dcd808fc",
          2846 => x"050c8053",
          2847 => x"81dcd808",
          2848 => x"8c050852",
          2849 => x"81dcd808",
          2850 => x"88050851",
          2851 => x"81df3f81",
          2852 => x"dccc0870",
          2853 => x"81dcd808",
          2854 => x"f8050c54",
          2855 => x"81dcd808",
          2856 => x"fc050880",
          2857 => x"2e903881",
          2858 => x"dcd808f8",
          2859 => x"05083081",
          2860 => x"dcd808f8",
          2861 => x"050c81dc",
          2862 => x"d808f805",
          2863 => x"087081dc",
          2864 => x"cc0c5489",
          2865 => x"3d0d81dc",
          2866 => x"d80c0481",
          2867 => x"dcd80802",
          2868 => x"81dcd80c",
          2869 => x"fb3d0d80",
          2870 => x"0b81dcd8",
          2871 => x"08fc050c",
          2872 => x"81dcd808",
          2873 => x"88050880",
          2874 => x"25993881",
          2875 => x"dcd80888",
          2876 => x"05083081",
          2877 => x"dcd80888",
          2878 => x"050c810b",
          2879 => x"81dcd808",
          2880 => x"fc050c81",
          2881 => x"dcd8088c",
          2882 => x"05088025",
          2883 => x"903881dc",
          2884 => x"d8088c05",
          2885 => x"083081dc",
          2886 => x"d8088c05",
          2887 => x"0c815381",
          2888 => x"dcd8088c",
          2889 => x"05085281",
          2890 => x"dcd80888",
          2891 => x"050851bd",
          2892 => x"3f81dccc",
          2893 => x"087081dc",
          2894 => x"d808f805",
          2895 => x"0c5481dc",
          2896 => x"d808fc05",
          2897 => x"08802e90",
          2898 => x"3881dcd8",
          2899 => x"08f80508",
          2900 => x"3081dcd8",
          2901 => x"08f8050c",
          2902 => x"81dcd808",
          2903 => x"f8050870",
          2904 => x"81dccc0c",
          2905 => x"54873d0d",
          2906 => x"81dcd80c",
          2907 => x"0481dcd8",
          2908 => x"080281dc",
          2909 => x"d80cfd3d",
          2910 => x"0d810b81",
          2911 => x"dcd808fc",
          2912 => x"050c800b",
          2913 => x"81dcd808",
          2914 => x"f8050c81",
          2915 => x"dcd8088c",
          2916 => x"050881dc",
          2917 => x"d8088805",
          2918 => x"0827b938",
          2919 => x"81dcd808",
          2920 => x"fc050880",
          2921 => x"2eae3880",
          2922 => x"0b81dcd8",
          2923 => x"088c0508",
          2924 => x"24a23881",
          2925 => x"dcd8088c",
          2926 => x"05081081",
          2927 => x"dcd8088c",
          2928 => x"050c81dc",
          2929 => x"d808fc05",
          2930 => x"081081dc",
          2931 => x"d808fc05",
          2932 => x"0cffb839",
          2933 => x"81dcd808",
          2934 => x"fc050880",
          2935 => x"2e80e138",
          2936 => x"81dcd808",
          2937 => x"8c050881",
          2938 => x"dcd80888",
          2939 => x"050826ad",
          2940 => x"3881dcd8",
          2941 => x"08880508",
          2942 => x"81dcd808",
          2943 => x"8c050831",
          2944 => x"81dcd808",
          2945 => x"88050c81",
          2946 => x"dcd808f8",
          2947 => x"050881dc",
          2948 => x"d808fc05",
          2949 => x"080781dc",
          2950 => x"d808f805",
          2951 => x"0c81dcd8",
          2952 => x"08fc0508",
          2953 => x"812a81dc",
          2954 => x"d808fc05",
          2955 => x"0c81dcd8",
          2956 => x"088c0508",
          2957 => x"812a81dc",
          2958 => x"d8088c05",
          2959 => x"0cff9539",
          2960 => x"81dcd808",
          2961 => x"90050880",
          2962 => x"2e933881",
          2963 => x"dcd80888",
          2964 => x"05087081",
          2965 => x"dcd808f4",
          2966 => x"050c5191",
          2967 => x"3981dcd8",
          2968 => x"08f80508",
          2969 => x"7081dcd8",
          2970 => x"08f4050c",
          2971 => x"5181dcd8",
          2972 => x"08f40508",
          2973 => x"81dccc0c",
          2974 => x"853d0d81",
          2975 => x"dcd80c04",
          2976 => x"fc3d0d76",
          2977 => x"7971028c",
          2978 => x"059f0533",
          2979 => x"57555355",
          2980 => x"8372278a",
          2981 => x"38748306",
          2982 => x"5170802e",
          2983 => x"a438ff12",
          2984 => x"5271ff2e",
          2985 => x"93387373",
          2986 => x"70810555",
          2987 => x"34ff1252",
          2988 => x"71ff2e09",
          2989 => x"8106ef38",
          2990 => x"7481dccc",
          2991 => x"0c863d0d",
          2992 => x"04747488",
          2993 => x"2b750770",
          2994 => x"71902b07",
          2995 => x"5154518f",
          2996 => x"7227a538",
          2997 => x"72717084",
          2998 => x"05530c72",
          2999 => x"71708405",
          3000 => x"530c7271",
          3001 => x"70840553",
          3002 => x"0c727170",
          3003 => x"8405530c",
          3004 => x"f0125271",
          3005 => x"8f26dd38",
          3006 => x"83722790",
          3007 => x"38727170",
          3008 => x"8405530c",
          3009 => x"fc125271",
          3010 => x"8326f238",
          3011 => x"7053ff8e",
          3012 => x"39fb3d0d",
          3013 => x"77797072",
          3014 => x"07830653",
          3015 => x"54527093",
          3016 => x"38717373",
          3017 => x"08545654",
          3018 => x"7173082e",
          3019 => x"80c63873",
          3020 => x"75545271",
          3021 => x"337081ff",
          3022 => x"06525470",
          3023 => x"802e9d38",
          3024 => x"72335570",
          3025 => x"752e0981",
          3026 => x"06953881",
          3027 => x"12811471",
          3028 => x"337081ff",
          3029 => x"06545654",
          3030 => x"5270e538",
          3031 => x"72335573",
          3032 => x"81ff0675",
          3033 => x"81ff0671",
          3034 => x"713181dc",
          3035 => x"cc0c5252",
          3036 => x"873d0d04",
          3037 => x"710970f7",
          3038 => x"fbfdff14",
          3039 => x"0670f884",
          3040 => x"82818006",
          3041 => x"51515170",
          3042 => x"97388414",
          3043 => x"84167108",
          3044 => x"54565471",
          3045 => x"75082edc",
          3046 => x"38737554",
          3047 => x"52ff9439",
          3048 => x"800b81dc",
          3049 => x"cc0c873d",
          3050 => x"0d04fe3d",
          3051 => x"0d805283",
          3052 => x"5371882b",
          3053 => x"5287863f",
          3054 => x"81dccc08",
          3055 => x"81ff0672",
          3056 => x"07ff1454",
          3057 => x"52728025",
          3058 => x"e8387181",
          3059 => x"dccc0c84",
          3060 => x"3d0d04fb",
          3061 => x"3d0d7770",
          3062 => x"08705353",
          3063 => x"5671802e",
          3064 => x"80ca3871",
          3065 => x"335170a0",
          3066 => x"2e098106",
          3067 => x"86388112",
          3068 => x"52f13971",
          3069 => x"53843981",
          3070 => x"13538073",
          3071 => x"337081ff",
          3072 => x"06535555",
          3073 => x"70a02e83",
          3074 => x"38815570",
          3075 => x"802e8438",
          3076 => x"74e53873",
          3077 => x"81ff0651",
          3078 => x"70a02e09",
          3079 => x"81068838",
          3080 => x"80737081",
          3081 => x"05553472",
          3082 => x"760c7151",
          3083 => x"7081dccc",
          3084 => x"0c873d0d",
          3085 => x"04fc3d0d",
          3086 => x"76537208",
          3087 => x"802e9138",
          3088 => x"863dfc05",
          3089 => x"5272519b",
          3090 => x"823f81dc",
          3091 => x"cc088538",
          3092 => x"80538339",
          3093 => x"74537281",
          3094 => x"dccc0c86",
          3095 => x"3d0d04fc",
          3096 => x"3d0d7682",
          3097 => x"1133ff05",
          3098 => x"52538152",
          3099 => x"708b2681",
          3100 => x"98388313",
          3101 => x"33ff0551",
          3102 => x"8252709e",
          3103 => x"26818a38",
          3104 => x"84133351",
          3105 => x"83527097",
          3106 => x"2680fe38",
          3107 => x"85133351",
          3108 => x"845270bb",
          3109 => x"2680f238",
          3110 => x"86133351",
          3111 => x"855270bb",
          3112 => x"2680e638",
          3113 => x"88132255",
          3114 => x"86527487",
          3115 => x"e72680d9",
          3116 => x"388a1322",
          3117 => x"54875273",
          3118 => x"87e72680",
          3119 => x"cc38810b",
          3120 => x"87c0989c",
          3121 => x"0c722287",
          3122 => x"c098bc0c",
          3123 => x"82133387",
          3124 => x"c098b80c",
          3125 => x"83133387",
          3126 => x"c098b40c",
          3127 => x"84133387",
          3128 => x"c098b00c",
          3129 => x"85133387",
          3130 => x"c098ac0c",
          3131 => x"86133387",
          3132 => x"c098a80c",
          3133 => x"7487c098",
          3134 => x"a40c7387",
          3135 => x"c098a00c",
          3136 => x"800b87c0",
          3137 => x"989c0c80",
          3138 => x"527181dc",
          3139 => x"cc0c863d",
          3140 => x"0d04f33d",
          3141 => x"0d7f5b87",
          3142 => x"c0989c5d",
          3143 => x"817d0c87",
          3144 => x"c098bc08",
          3145 => x"5e7d7b23",
          3146 => x"87c098b8",
          3147 => x"085a7982",
          3148 => x"1c3487c0",
          3149 => x"98b4085a",
          3150 => x"79831c34",
          3151 => x"87c098b0",
          3152 => x"085a7984",
          3153 => x"1c3487c0",
          3154 => x"98ac085a",
          3155 => x"79851c34",
          3156 => x"87c098a8",
          3157 => x"085a7986",
          3158 => x"1c3487c0",
          3159 => x"98a4085c",
          3160 => x"7b881c23",
          3161 => x"87c098a0",
          3162 => x"085a798a",
          3163 => x"1c23807d",
          3164 => x"0c7983ff",
          3165 => x"ff06597b",
          3166 => x"83ffff06",
          3167 => x"58861b33",
          3168 => x"57851b33",
          3169 => x"56841b33",
          3170 => x"55831b33",
          3171 => x"54821b33",
          3172 => x"537d83ff",
          3173 => x"ff065281",
          3174 => x"c5cc5194",
          3175 => x"c73f8f3d",
          3176 => x"0d04ff3d",
          3177 => x"0d028f05",
          3178 => x"33703070",
          3179 => x"9f2a5152",
          3180 => x"52700b0b",
          3181 => x"81d8f434",
          3182 => x"833d0d04",
          3183 => x"fb3d0d77",
          3184 => x"0b0b81d8",
          3185 => x"f4337081",
          3186 => x"ff065755",
          3187 => x"5687c094",
          3188 => x"84517480",
          3189 => x"2e863887",
          3190 => x"c0949451",
          3191 => x"70087096",
          3192 => x"2a708106",
          3193 => x"53545270",
          3194 => x"802e8c38",
          3195 => x"71912a70",
          3196 => x"81065151",
          3197 => x"70d73872",
          3198 => x"81327081",
          3199 => x"06515170",
          3200 => x"802e8d38",
          3201 => x"71932a70",
          3202 => x"81065151",
          3203 => x"70ffbe38",
          3204 => x"7381ff06",
          3205 => x"5187c094",
          3206 => x"80527080",
          3207 => x"2e863887",
          3208 => x"c0949052",
          3209 => x"75720c75",
          3210 => x"81dccc0c",
          3211 => x"873d0d04",
          3212 => x"fb3d0d02",
          3213 => x"9f05330b",
          3214 => x"0b81d8f4",
          3215 => x"337081ff",
          3216 => x"06575556",
          3217 => x"87c09484",
          3218 => x"5174802e",
          3219 => x"863887c0",
          3220 => x"94945170",
          3221 => x"0870962a",
          3222 => x"70810653",
          3223 => x"54527080",
          3224 => x"2e8c3871",
          3225 => x"912a7081",
          3226 => x"06515170",
          3227 => x"d7387281",
          3228 => x"32708106",
          3229 => x"51517080",
          3230 => x"2e8d3871",
          3231 => x"932a7081",
          3232 => x"06515170",
          3233 => x"ffbe3873",
          3234 => x"81ff0651",
          3235 => x"87c09480",
          3236 => x"5270802e",
          3237 => x"863887c0",
          3238 => x"94905275",
          3239 => x"720c873d",
          3240 => x"0d04f93d",
          3241 => x"0d795480",
          3242 => x"74337081",
          3243 => x"ff065353",
          3244 => x"5770772e",
          3245 => x"80fe3871",
          3246 => x"81ff0681",
          3247 => x"150b0b81",
          3248 => x"d8f43370",
          3249 => x"81ff0659",
          3250 => x"57555887",
          3251 => x"c0948451",
          3252 => x"75802e86",
          3253 => x"3887c094",
          3254 => x"94517008",
          3255 => x"70962a70",
          3256 => x"81065354",
          3257 => x"5270802e",
          3258 => x"8c387191",
          3259 => x"2a708106",
          3260 => x"515170d7",
          3261 => x"38728132",
          3262 => x"70810651",
          3263 => x"5170802e",
          3264 => x"8d387193",
          3265 => x"2a708106",
          3266 => x"515170ff",
          3267 => x"be387481",
          3268 => x"ff065187",
          3269 => x"c0948052",
          3270 => x"70802e86",
          3271 => x"3887c094",
          3272 => x"90527772",
          3273 => x"0c811774",
          3274 => x"337081ff",
          3275 => x"06535357",
          3276 => x"70ff8438",
          3277 => x"7681dccc",
          3278 => x"0c893d0d",
          3279 => x"04fe3d0d",
          3280 => x"0b0b81d8",
          3281 => x"f4337081",
          3282 => x"ff065452",
          3283 => x"87c09484",
          3284 => x"5172802e",
          3285 => x"863887c0",
          3286 => x"94945170",
          3287 => x"0870822a",
          3288 => x"70810651",
          3289 => x"51517080",
          3290 => x"2ee23871",
          3291 => x"81ff0651",
          3292 => x"87c09480",
          3293 => x"5270802e",
          3294 => x"863887c0",
          3295 => x"94905271",
          3296 => x"087081ff",
          3297 => x"0681dccc",
          3298 => x"0c51843d",
          3299 => x"0d04fe3d",
          3300 => x"0d0b0b81",
          3301 => x"d8f43370",
          3302 => x"81ff0652",
          3303 => x"5387c094",
          3304 => x"84527080",
          3305 => x"2e863887",
          3306 => x"c0949452",
          3307 => x"71087082",
          3308 => x"2a708106",
          3309 => x"515151ff",
          3310 => x"5270802e",
          3311 => x"a0387281",
          3312 => x"ff065187",
          3313 => x"c0948052",
          3314 => x"70802e86",
          3315 => x"3887c094",
          3316 => x"90527108",
          3317 => x"70982b70",
          3318 => x"982c5153",
          3319 => x"517181dc",
          3320 => x"cc0c843d",
          3321 => x"0d04ff3d",
          3322 => x"0d87c09e",
          3323 => x"8008709c",
          3324 => x"2a8a0651",
          3325 => x"5170802e",
          3326 => x"84b43887",
          3327 => x"c09ea408",
          3328 => x"81d8f80c",
          3329 => x"87c09ea8",
          3330 => x"0881d8fc",
          3331 => x"0c87c09e",
          3332 => x"940881d9",
          3333 => x"800c87c0",
          3334 => x"9e980881",
          3335 => x"d9840c87",
          3336 => x"c09e9c08",
          3337 => x"81d9880c",
          3338 => x"87c09ea0",
          3339 => x"0881d98c",
          3340 => x"0c87c09e",
          3341 => x"ac0881d9",
          3342 => x"900c87c0",
          3343 => x"9eb00881",
          3344 => x"d9940c87",
          3345 => x"c09eb408",
          3346 => x"81d9980c",
          3347 => x"87c09eb8",
          3348 => x"0881d99c",
          3349 => x"0c87c09e",
          3350 => x"bc0881d9",
          3351 => x"a00c87c0",
          3352 => x"9ec00881",
          3353 => x"d9a40c87",
          3354 => x"c09ec408",
          3355 => x"81d9a80c",
          3356 => x"87c09e80",
          3357 => x"08517081",
          3358 => x"d9ac2387",
          3359 => x"c09e8408",
          3360 => x"81d9b00c",
          3361 => x"87c09e88",
          3362 => x"0881d9b4",
          3363 => x"0c87c09e",
          3364 => x"8c0881d9",
          3365 => x"b80c810b",
          3366 => x"81d9bc34",
          3367 => x"800b87c0",
          3368 => x"9e900870",
          3369 => x"84800a06",
          3370 => x"51525270",
          3371 => x"802e8338",
          3372 => x"81527181",
          3373 => x"d9bd3480",
          3374 => x"0b87c09e",
          3375 => x"90087088",
          3376 => x"800a0651",
          3377 => x"52527080",
          3378 => x"2e833881",
          3379 => x"527181d9",
          3380 => x"be34800b",
          3381 => x"87c09e90",
          3382 => x"08709080",
          3383 => x"0a065152",
          3384 => x"5270802e",
          3385 => x"83388152",
          3386 => x"7181d9bf",
          3387 => x"34800b87",
          3388 => x"c09e9008",
          3389 => x"70888080",
          3390 => x"06515252",
          3391 => x"70802e83",
          3392 => x"38815271",
          3393 => x"81d9c034",
          3394 => x"800b87c0",
          3395 => x"9e900870",
          3396 => x"a0808006",
          3397 => x"51525270",
          3398 => x"802e8338",
          3399 => x"81527181",
          3400 => x"d9c13480",
          3401 => x"0b87c09e",
          3402 => x"90087090",
          3403 => x"80800651",
          3404 => x"52527080",
          3405 => x"2e833881",
          3406 => x"527181d9",
          3407 => x"c234800b",
          3408 => x"87c09e90",
          3409 => x"08708480",
          3410 => x"80065152",
          3411 => x"5270802e",
          3412 => x"83388152",
          3413 => x"7181d9c3",
          3414 => x"34800b87",
          3415 => x"c09e9008",
          3416 => x"70828080",
          3417 => x"06515252",
          3418 => x"70802e83",
          3419 => x"38815271",
          3420 => x"81d9c434",
          3421 => x"800b87c0",
          3422 => x"9e900870",
          3423 => x"81808006",
          3424 => x"51525270",
          3425 => x"802e8338",
          3426 => x"81527181",
          3427 => x"d9c53480",
          3428 => x"0b87c09e",
          3429 => x"90087080",
          3430 => x"c0800651",
          3431 => x"52527080",
          3432 => x"2e833881",
          3433 => x"527181d9",
          3434 => x"c634800b",
          3435 => x"87c09e90",
          3436 => x"0870a080",
          3437 => x"06515252",
          3438 => x"70802e83",
          3439 => x"38815271",
          3440 => x"81d9c734",
          3441 => x"87c09e90",
          3442 => x"08709880",
          3443 => x"06708a2a",
          3444 => x"51515170",
          3445 => x"81d9c834",
          3446 => x"800b87c0",
          3447 => x"9e900870",
          3448 => x"84800651",
          3449 => x"52527080",
          3450 => x"2e833881",
          3451 => x"527181d9",
          3452 => x"c93487c0",
          3453 => x"9e900870",
          3454 => x"83f00670",
          3455 => x"842a5151",
          3456 => x"517081d9",
          3457 => x"ca34800b",
          3458 => x"87c09e90",
          3459 => x"08708806",
          3460 => x"51525270",
          3461 => x"802e8338",
          3462 => x"81527181",
          3463 => x"d9cb3487",
          3464 => x"c09e9008",
          3465 => x"70870651",
          3466 => x"517081d9",
          3467 => x"cc34833d",
          3468 => x"0d04fb3d",
          3469 => x"0d81c5e4",
          3470 => x"5185c53f",
          3471 => x"81d9bc33",
          3472 => x"5473802e",
          3473 => x"883881c5",
          3474 => x"f85185b4",
          3475 => x"3f81c68c",
          3476 => x"5185ad3f",
          3477 => x"81d9be33",
          3478 => x"5473802e",
          3479 => x"933881d9",
          3480 => x"980881d9",
          3481 => x"9c081154",
          3482 => x"5281c6a4",
          3483 => x"518af53f",
          3484 => x"81d9c333",
          3485 => x"5473802e",
          3486 => x"933881d9",
          3487 => x"900881d9",
          3488 => x"94081154",
          3489 => x"5281c6c0",
          3490 => x"518ad93f",
          3491 => x"81d9c033",
          3492 => x"5473802e",
          3493 => x"933881d8",
          3494 => x"f80881d8",
          3495 => x"fc081154",
          3496 => x"5281c6dc",
          3497 => x"518abd3f",
          3498 => x"81d9c133",
          3499 => x"5473802e",
          3500 => x"933881d9",
          3501 => x"800881d9",
          3502 => x"84081154",
          3503 => x"5281c6f8",
          3504 => x"518aa13f",
          3505 => x"81d9c233",
          3506 => x"5473802e",
          3507 => x"933881d9",
          3508 => x"880881d9",
          3509 => x"8c081154",
          3510 => x"5281c794",
          3511 => x"518a853f",
          3512 => x"81d9c733",
          3513 => x"5473802e",
          3514 => x"8d3881d9",
          3515 => x"c8335281",
          3516 => x"c7b05189",
          3517 => x"ef3f81d9",
          3518 => x"cb335473",
          3519 => x"802e8d38",
          3520 => x"81d9cc33",
          3521 => x"5281c7d0",
          3522 => x"5189d93f",
          3523 => x"81d9c933",
          3524 => x"5473802e",
          3525 => x"8d3881d9",
          3526 => x"ca335281",
          3527 => x"c7f05189",
          3528 => x"c33f81d9",
          3529 => x"bd335473",
          3530 => x"802e8838",
          3531 => x"81c89051",
          3532 => x"83ce3f81",
          3533 => x"d9bf3354",
          3534 => x"73802e88",
          3535 => x"3881c8a4",
          3536 => x"5183bd3f",
          3537 => x"81d9c433",
          3538 => x"5473802e",
          3539 => x"883881c8",
          3540 => x"b05183ac",
          3541 => x"3f81d9c5",
          3542 => x"33547380",
          3543 => x"2e883881",
          3544 => x"c8bc5183",
          3545 => x"9b3f81d9",
          3546 => x"c6335473",
          3547 => x"802e8838",
          3548 => x"81c8c851",
          3549 => x"838a3f81",
          3550 => x"c8d45183",
          3551 => x"833f81d9",
          3552 => x"a0085281",
          3553 => x"c8e05188",
          3554 => x"db3f81d9",
          3555 => x"a4085281",
          3556 => x"c9885188",
          3557 => x"cf3f81d9",
          3558 => x"a8085281",
          3559 => x"c9b05188",
          3560 => x"c33f81c9",
          3561 => x"d85182d8",
          3562 => x"3f81d9ac",
          3563 => x"225281c9",
          3564 => x"e05188b0",
          3565 => x"3f81d9b0",
          3566 => x"0856bd84",
          3567 => x"c0527551",
          3568 => x"e7b73f81",
          3569 => x"dccc08bd",
          3570 => x"84c02976",
          3571 => x"71315454",
          3572 => x"81dccc08",
          3573 => x"5281ca88",
          3574 => x"5188893f",
          3575 => x"81d9c333",
          3576 => x"5473802e",
          3577 => x"a83881d9",
          3578 => x"b40856bd",
          3579 => x"84c05275",
          3580 => x"51e7863f",
          3581 => x"81dccc08",
          3582 => x"bd84c029",
          3583 => x"76713154",
          3584 => x"5481dccc",
          3585 => x"085281ca",
          3586 => x"b45187d8",
          3587 => x"3f81d9be",
          3588 => x"33547380",
          3589 => x"2ea83881",
          3590 => x"d9b80856",
          3591 => x"bd84c052",
          3592 => x"7551e6d5",
          3593 => x"3f81dccc",
          3594 => x"08bd84c0",
          3595 => x"29767131",
          3596 => x"545481dc",
          3597 => x"cc085281",
          3598 => x"cae05187",
          3599 => x"a73f81d6",
          3600 => x"c45181bc",
          3601 => x"3f873d0d",
          3602 => x"04fe3d0d",
          3603 => x"02920533",
          3604 => x"ff055271",
          3605 => x"8426aa38",
          3606 => x"71842981",
          3607 => x"c4e80552",
          3608 => x"71080481",
          3609 => x"cb8c519d",
          3610 => x"3981cb94",
          3611 => x"51973981",
          3612 => x"cb9c5191",
          3613 => x"3981cba4",
          3614 => x"518b3981",
          3615 => x"cba85185",
          3616 => x"3981cbb0",
          3617 => x"5180f93f",
          3618 => x"843d0d04",
          3619 => x"7188800c",
          3620 => x"04800b87",
          3621 => x"c096840c",
          3622 => x"0481d9d0",
          3623 => x"0887c096",
          3624 => x"840c04fe",
          3625 => x"3d0d0293",
          3626 => x"05335372",
          3627 => x"8a2e0981",
          3628 => x"0685388d",
          3629 => x"51ed3f81",
          3630 => x"dce40852",
          3631 => x"71802e90",
          3632 => x"38727234",
          3633 => x"81dce408",
          3634 => x"810581dc",
          3635 => x"e40c8f39",
          3636 => x"81dcdc08",
          3637 => x"5271802e",
          3638 => x"85387251",
          3639 => x"712d843d",
          3640 => x"0d04fe3d",
          3641 => x"0d029705",
          3642 => x"3381dcdc",
          3643 => x"087681dc",
          3644 => x"dc0c5451",
          3645 => x"ffad3f72",
          3646 => x"81dcdc0c",
          3647 => x"843d0d04",
          3648 => x"fd3d0d75",
          3649 => x"54733370",
          3650 => x"81ff0653",
          3651 => x"5371802e",
          3652 => x"8e387281",
          3653 => x"ff065181",
          3654 => x"1454ff87",
          3655 => x"3fe73985",
          3656 => x"3d0d04fc",
          3657 => x"3d0d7781",
          3658 => x"dcdc0878",
          3659 => x"81dcdc0c",
          3660 => x"56547333",
          3661 => x"7081ff06",
          3662 => x"53537180",
          3663 => x"2e8e3872",
          3664 => x"81ff0651",
          3665 => x"811454fe",
          3666 => x"da3fe739",
          3667 => x"7481dcdc",
          3668 => x"0c863d0d",
          3669 => x"04ec3d0d",
          3670 => x"66685959",
          3671 => x"78708105",
          3672 => x"5a335675",
          3673 => x"802e84f8",
          3674 => x"3875a52e",
          3675 => x"09810682",
          3676 => x"de388070",
          3677 => x"7a708105",
          3678 => x"5c33585b",
          3679 => x"5b75b02e",
          3680 => x"09810685",
          3681 => x"38815a8b",
          3682 => x"3975ad2e",
          3683 => x"0981068a",
          3684 => x"38825a78",
          3685 => x"7081055a",
          3686 => x"335675aa",
          3687 => x"2e098106",
          3688 => x"92387784",
          3689 => x"1971087b",
          3690 => x"7081055d",
          3691 => x"33595d59",
          3692 => x"539d39d0",
          3693 => x"16537289",
          3694 => x"2695387a",
          3695 => x"88297b10",
          3696 => x"057605d0",
          3697 => x"05797081",
          3698 => x"055b3357",
          3699 => x"5be53975",
          3700 => x"80ec3270",
          3701 => x"30707207",
          3702 => x"80257880",
          3703 => x"cc327030",
          3704 => x"70720780",
          3705 => x"25730753",
          3706 => x"54585155",
          3707 => x"5373802e",
          3708 => x"8c387984",
          3709 => x"07797081",
          3710 => x"055b3357",
          3711 => x"5a75802e",
          3712 => x"83de3875",
          3713 => x"5480e076",
          3714 => x"278938e0",
          3715 => x"167081ff",
          3716 => x"06555373",
          3717 => x"80cf2e81",
          3718 => x"aa387380",
          3719 => x"cf24a238",
          3720 => x"7380c32e",
          3721 => x"818e3873",
          3722 => x"80c3248b",
          3723 => x"387380c2",
          3724 => x"2e818c38",
          3725 => x"81993973",
          3726 => x"80c42e81",
          3727 => x"8a38818f",
          3728 => x"397380d5",
          3729 => x"2e818038",
          3730 => x"7380d524",
          3731 => x"8a387380",
          3732 => x"d32e8e38",
          3733 => x"80f93973",
          3734 => x"80d82e80",
          3735 => x"ee3880ef",
          3736 => x"39778419",
          3737 => x"71085659",
          3738 => x"53807433",
          3739 => x"54557275",
          3740 => x"2e8d3881",
          3741 => x"15701570",
          3742 => x"33515455",
          3743 => x"72f53879",
          3744 => x"812a5690",
          3745 => x"39748116",
          3746 => x"5653727b",
          3747 => x"278f38a0",
          3748 => x"51fc903f",
          3749 => x"75810653",
          3750 => x"72802ee9",
          3751 => x"387351fc",
          3752 => x"df3f7481",
          3753 => x"16565372",
          3754 => x"7b27fdb0",
          3755 => x"38a051fb",
          3756 => x"f23fef39",
          3757 => x"77841983",
          3758 => x"12335359",
          3759 => x"53933982",
          3760 => x"5c953988",
          3761 => x"5c91398a",
          3762 => x"5c8d3990",
          3763 => x"5c893975",
          3764 => x"51fbd03f",
          3765 => x"fd863979",
          3766 => x"822a7081",
          3767 => x"06515372",
          3768 => x"802e8838",
          3769 => x"77841959",
          3770 => x"53863984",
          3771 => x"18785458",
          3772 => x"72087480",
          3773 => x"c4327030",
          3774 => x"70720780",
          3775 => x"25515555",
          3776 => x"55748025",
          3777 => x"8d387280",
          3778 => x"2e883874",
          3779 => x"307a9007",
          3780 => x"5b55800b",
          3781 => x"8f3d5e57",
          3782 => x"7b527451",
          3783 => x"e18e3f81",
          3784 => x"dccc0881",
          3785 => x"ff067c53",
          3786 => x"755254e0",
          3787 => x"cc3f81dc",
          3788 => x"cc085589",
          3789 => x"74279238",
          3790 => x"a7145375",
          3791 => x"80f82e84",
          3792 => x"38871453",
          3793 => x"7281ff06",
          3794 => x"54b01453",
          3795 => x"727d7081",
          3796 => x"055f3481",
          3797 => x"17753070",
          3798 => x"77079f2a",
          3799 => x"51545776",
          3800 => x"9f268538",
          3801 => x"72ffb138",
          3802 => x"79842a70",
          3803 => x"81065153",
          3804 => x"72802e8e",
          3805 => x"38963d77",
          3806 => x"05e00553",
          3807 => x"ad733481",
          3808 => x"1757767a",
          3809 => x"81065455",
          3810 => x"b0547283",
          3811 => x"38a05479",
          3812 => x"812a7081",
          3813 => x"06545672",
          3814 => x"9f388117",
          3815 => x"55767b27",
          3816 => x"97387351",
          3817 => x"f9fd3f75",
          3818 => x"81065372",
          3819 => x"8b387481",
          3820 => x"1656537a",
          3821 => x"7326eb38",
          3822 => x"963d7705",
          3823 => x"e00553ff",
          3824 => x"17ff1470",
          3825 => x"33535457",
          3826 => x"f9d93f76",
          3827 => x"f2387481",
          3828 => x"16565372",
          3829 => x"7b27fb84",
          3830 => x"38a051f9",
          3831 => x"c63fef39",
          3832 => x"963d0d04",
          3833 => x"fd3d0d86",
          3834 => x"3d707084",
          3835 => x"05520855",
          3836 => x"527351fa",
          3837 => x"e03f853d",
          3838 => x"0d04fe3d",
          3839 => x"0d7481dc",
          3840 => x"e40c853d",
          3841 => x"88055275",
          3842 => x"51faca3f",
          3843 => x"81dce408",
          3844 => x"53807334",
          3845 => x"800b81dc",
          3846 => x"e40c843d",
          3847 => x"0d04fd3d",
          3848 => x"0d81dcdc",
          3849 => x"087681dc",
          3850 => x"dc0c873d",
          3851 => x"88055377",
          3852 => x"5253faa1",
          3853 => x"3f7281dc",
          3854 => x"dc0c853d",
          3855 => x"0d04fb3d",
          3856 => x"0d777981",
          3857 => x"dce00870",
          3858 => x"56545755",
          3859 => x"80547180",
          3860 => x"2e80e038",
          3861 => x"81dce008",
          3862 => x"52712d81",
          3863 => x"dccc0881",
          3864 => x"ff065372",
          3865 => x"802e80cb",
          3866 => x"38728d2e",
          3867 => x"b9387288",
          3868 => x"32703070",
          3869 => x"80255151",
          3870 => x"5273802e",
          3871 => x"8b387180",
          3872 => x"2e8638ff",
          3873 => x"14549739",
          3874 => x"9f7325c8",
          3875 => x"38ff1652",
          3876 => x"737225c0",
          3877 => x"38741452",
          3878 => x"72723481",
          3879 => x"14547251",
          3880 => x"f8813fff",
          3881 => x"af397315",
          3882 => x"52807234",
          3883 => x"8a51f7f3",
          3884 => x"3f815372",
          3885 => x"81dccc0c",
          3886 => x"873d0d04",
          3887 => x"fe3d0d81",
          3888 => x"dce00875",
          3889 => x"81dce00c",
          3890 => x"77537652",
          3891 => x"53feef3f",
          3892 => x"7281dce0",
          3893 => x"0c843d0d",
          3894 => x"04f83d0d",
          3895 => x"7a7c5a56",
          3896 => x"80707a0c",
          3897 => x"58750870",
          3898 => x"33555373",
          3899 => x"a02e0981",
          3900 => x"06873881",
          3901 => x"13760ced",
          3902 => x"3973ad2e",
          3903 => x"0981068e",
          3904 => x"38817608",
          3905 => x"11770c76",
          3906 => x"08703356",
          3907 => x"545873b0",
          3908 => x"2e098106",
          3909 => x"80c23875",
          3910 => x"08810576",
          3911 => x"0c750870",
          3912 => x"33555373",
          3913 => x"80e22e8b",
          3914 => x"38905773",
          3915 => x"80f82e85",
          3916 => x"388f3982",
          3917 => x"57811376",
          3918 => x"0c750870",
          3919 => x"335553ac",
          3920 => x"398155a0",
          3921 => x"742780fa",
          3922 => x"38d01453",
          3923 => x"80558857",
          3924 => x"89732798",
          3925 => x"3880eb39",
          3926 => x"d0145380",
          3927 => x"55728926",
          3928 => x"80e03886",
          3929 => x"39805580",
          3930 => x"d9398a57",
          3931 => x"8055a074",
          3932 => x"2780c238",
          3933 => x"80e07427",
          3934 => x"8938e014",
          3935 => x"7081ff06",
          3936 => x"5553d014",
          3937 => x"7081ff06",
          3938 => x"55539074",
          3939 => x"278e38f9",
          3940 => x"147081ff",
          3941 => x"06555389",
          3942 => x"7427ca38",
          3943 => x"737727c5",
          3944 => x"38747729",
          3945 => x"14760881",
          3946 => x"05770c76",
          3947 => x"08703356",
          3948 => x"5455ffba",
          3949 => x"3977802e",
          3950 => x"84387430",
          3951 => x"5574790c",
          3952 => x"81557481",
          3953 => x"dccc0c8a",
          3954 => x"3d0d04f8",
          3955 => x"3d0d7a7c",
          3956 => x"5a568070",
          3957 => x"7a0c5875",
          3958 => x"08703355",
          3959 => x"5373a02e",
          3960 => x"09810687",
          3961 => x"38811376",
          3962 => x"0ced3973",
          3963 => x"ad2e0981",
          3964 => x"068e3881",
          3965 => x"76081177",
          3966 => x"0c760870",
          3967 => x"33565458",
          3968 => x"73b02e09",
          3969 => x"810680c2",
          3970 => x"38750881",
          3971 => x"05760c75",
          3972 => x"08703355",
          3973 => x"537380e2",
          3974 => x"2e8b3890",
          3975 => x"577380f8",
          3976 => x"2e85388f",
          3977 => x"39825781",
          3978 => x"13760c75",
          3979 => x"08703355",
          3980 => x"53ac3981",
          3981 => x"55a07427",
          3982 => x"80fa38d0",
          3983 => x"14538055",
          3984 => x"88578973",
          3985 => x"27983880",
          3986 => x"eb39d014",
          3987 => x"53805572",
          3988 => x"892680e0",
          3989 => x"38863980",
          3990 => x"5580d939",
          3991 => x"8a578055",
          3992 => x"a0742780",
          3993 => x"c23880e0",
          3994 => x"74278938",
          3995 => x"e0147081",
          3996 => x"ff065553",
          3997 => x"d0147081",
          3998 => x"ff065553",
          3999 => x"9074278e",
          4000 => x"38f91470",
          4001 => x"81ff0655",
          4002 => x"53897427",
          4003 => x"ca387377",
          4004 => x"27c53874",
          4005 => x"77291476",
          4006 => x"08810577",
          4007 => x"0c760870",
          4008 => x"33565455",
          4009 => x"ffba3977",
          4010 => x"802e8438",
          4011 => x"74305574",
          4012 => x"790c8155",
          4013 => x"7481dccc",
          4014 => x"0c8a3d0d",
          4015 => x"04ff3d0d",
          4016 => x"028f0533",
          4017 => x"51815270",
          4018 => x"72268738",
          4019 => x"81d9d411",
          4020 => x"33527181",
          4021 => x"dccc0c83",
          4022 => x"3d0d04fc",
          4023 => x"3d0d029b",
          4024 => x"05330284",
          4025 => x"059f0533",
          4026 => x"56538351",
          4027 => x"72812680",
          4028 => x"e0387284",
          4029 => x"2b87c092",
          4030 => x"8c115351",
          4031 => x"88547480",
          4032 => x"2e843881",
          4033 => x"88547372",
          4034 => x"0c87c092",
          4035 => x"8c115181",
          4036 => x"710c850b",
          4037 => x"87c0988c",
          4038 => x"0c705271",
          4039 => x"08708206",
          4040 => x"51517080",
          4041 => x"2e8a3887",
          4042 => x"c0988c08",
          4043 => x"5170ec38",
          4044 => x"7108fc80",
          4045 => x"80065271",
          4046 => x"923887c0",
          4047 => x"988c0851",
          4048 => x"70802e87",
          4049 => x"387181d9",
          4050 => x"d4143481",
          4051 => x"d9d41333",
          4052 => x"517081dc",
          4053 => x"cc0c863d",
          4054 => x"0d04f33d",
          4055 => x"0d606264",
          4056 => x"028c05bf",
          4057 => x"05335740",
          4058 => x"585b8374",
          4059 => x"525afecd",
          4060 => x"3f81dccc",
          4061 => x"0881067a",
          4062 => x"54527181",
          4063 => x"be387172",
          4064 => x"75842b87",
          4065 => x"c0928011",
          4066 => x"87c0928c",
          4067 => x"1287c092",
          4068 => x"8413415a",
          4069 => x"40575a58",
          4070 => x"850b87c0",
          4071 => x"988c0c76",
          4072 => x"7d0c8476",
          4073 => x"0c750870",
          4074 => x"852a7081",
          4075 => x"06515354",
          4076 => x"71802e8e",
          4077 => x"387b0852",
          4078 => x"717b7081",
          4079 => x"055d3481",
          4080 => x"19598074",
          4081 => x"a2065353",
          4082 => x"71732e83",
          4083 => x"38815378",
          4084 => x"83ff268f",
          4085 => x"3872802e",
          4086 => x"8a3887c0",
          4087 => x"988c0852",
          4088 => x"71c33887",
          4089 => x"c0988c08",
          4090 => x"5271802e",
          4091 => x"87387884",
          4092 => x"802e9938",
          4093 => x"81760c87",
          4094 => x"c0928c15",
          4095 => x"53720870",
          4096 => x"82065152",
          4097 => x"71f738ff",
          4098 => x"1a5a8d39",
          4099 => x"84801781",
          4100 => x"197081ff",
          4101 => x"065a5357",
          4102 => x"79802e90",
          4103 => x"3873fc80",
          4104 => x"80065271",
          4105 => x"87387d78",
          4106 => x"26feed38",
          4107 => x"73fc8080",
          4108 => x"06527180",
          4109 => x"2e833881",
          4110 => x"52715372",
          4111 => x"81dccc0c",
          4112 => x"8f3d0d04",
          4113 => x"f33d0d60",
          4114 => x"6264028c",
          4115 => x"05bf0533",
          4116 => x"5740585b",
          4117 => x"83598074",
          4118 => x"5258fce1",
          4119 => x"3f81dccc",
          4120 => x"08810679",
          4121 => x"54527178",
          4122 => x"2e098106",
          4123 => x"81b13877",
          4124 => x"74842b87",
          4125 => x"c0928011",
          4126 => x"87c0928c",
          4127 => x"1287c092",
          4128 => x"84134059",
          4129 => x"5f565a85",
          4130 => x"0b87c098",
          4131 => x"8c0c767d",
          4132 => x"0c82760c",
          4133 => x"80587508",
          4134 => x"70842a70",
          4135 => x"81065153",
          4136 => x"5471802e",
          4137 => x"8c387a70",
          4138 => x"81055c33",
          4139 => x"7c0c8118",
          4140 => x"5873812a",
          4141 => x"70810651",
          4142 => x"5271802e",
          4143 => x"8a3887c0",
          4144 => x"988c0852",
          4145 => x"71d03887",
          4146 => x"c0988c08",
          4147 => x"5271802e",
          4148 => x"87387784",
          4149 => x"802e9938",
          4150 => x"81760c87",
          4151 => x"c0928c15",
          4152 => x"53720870",
          4153 => x"82065152",
          4154 => x"71f738ff",
          4155 => x"19598d39",
          4156 => x"811a7081",
          4157 => x"ff068480",
          4158 => x"19595b52",
          4159 => x"78802e90",
          4160 => x"3873fc80",
          4161 => x"80065271",
          4162 => x"87387d7a",
          4163 => x"26fef838",
          4164 => x"73fc8080",
          4165 => x"06527180",
          4166 => x"2e833881",
          4167 => x"52715372",
          4168 => x"81dccc0c",
          4169 => x"8f3d0d04",
          4170 => x"fa3d0d7a",
          4171 => x"028405a3",
          4172 => x"05330288",
          4173 => x"05a70533",
          4174 => x"71545456",
          4175 => x"57fafe3f",
          4176 => x"81dccc08",
          4177 => x"81065383",
          4178 => x"547280fe",
          4179 => x"38850b87",
          4180 => x"c0988c0c",
          4181 => x"81567176",
          4182 => x"2e80dc38",
          4183 => x"71762493",
          4184 => x"3874842b",
          4185 => x"87c0928c",
          4186 => x"11545471",
          4187 => x"802e8d38",
          4188 => x"80d43971",
          4189 => x"832e80c6",
          4190 => x"3880cb39",
          4191 => x"72087081",
          4192 => x"2a708106",
          4193 => x"51515271",
          4194 => x"802e8a38",
          4195 => x"87c0988c",
          4196 => x"085271e8",
          4197 => x"3887c098",
          4198 => x"8c085271",
          4199 => x"96388173",
          4200 => x"0c87c092",
          4201 => x"8c145372",
          4202 => x"08708206",
          4203 => x"515271f7",
          4204 => x"38963980",
          4205 => x"56923988",
          4206 => x"800a770c",
          4207 => x"85398180",
          4208 => x"770c7256",
          4209 => x"83398456",
          4210 => x"75547381",
          4211 => x"dccc0c88",
          4212 => x"3d0d04fe",
          4213 => x"3d0d7481",
          4214 => x"11337133",
          4215 => x"71882b07",
          4216 => x"81dccc0c",
          4217 => x"5351843d",
          4218 => x"0d04fd3d",
          4219 => x"0d758311",
          4220 => x"33821233",
          4221 => x"71902b71",
          4222 => x"882b0781",
          4223 => x"14337072",
          4224 => x"07882b75",
          4225 => x"33710781",
          4226 => x"dccc0c52",
          4227 => x"53545654",
          4228 => x"52853d0d",
          4229 => x"04ff3d0d",
          4230 => x"73028405",
          4231 => x"92052252",
          4232 => x"52707270",
          4233 => x"81055434",
          4234 => x"70882a51",
          4235 => x"70723483",
          4236 => x"3d0d04ff",
          4237 => x"3d0d7375",
          4238 => x"52527072",
          4239 => x"70810554",
          4240 => x"3470882a",
          4241 => x"51707270",
          4242 => x"81055434",
          4243 => x"70882a51",
          4244 => x"70727081",
          4245 => x"05543470",
          4246 => x"882a5170",
          4247 => x"7234833d",
          4248 => x"0d04fe3d",
          4249 => x"0d767577",
          4250 => x"54545170",
          4251 => x"802e9238",
          4252 => x"71708105",
          4253 => x"53337370",
          4254 => x"81055534",
          4255 => x"ff1151eb",
          4256 => x"39843d0d",
          4257 => x"04fe3d0d",
          4258 => x"75777654",
          4259 => x"52537272",
          4260 => x"70810554",
          4261 => x"34ff1151",
          4262 => x"70f43884",
          4263 => x"3d0d04fc",
          4264 => x"3d0d7877",
          4265 => x"79565653",
          4266 => x"74708105",
          4267 => x"56337470",
          4268 => x"81055633",
          4269 => x"717131ff",
          4270 => x"16565252",
          4271 => x"5272802e",
          4272 => x"86387180",
          4273 => x"2ee23871",
          4274 => x"81dccc0c",
          4275 => x"863d0d04",
          4276 => x"fe3d0d74",
          4277 => x"76545189",
          4278 => x"3971732e",
          4279 => x"8a388111",
          4280 => x"51703352",
          4281 => x"71f33870",
          4282 => x"3381dccc",
          4283 => x"0c843d0d",
          4284 => x"04800b81",
          4285 => x"dccc0c04",
          4286 => x"800b81dc",
          4287 => x"cc0c04f7",
          4288 => x"3d0d7b56",
          4289 => x"800b8317",
          4290 => x"33565a74",
          4291 => x"7a2e80d6",
          4292 => x"388154b0",
          4293 => x"160853b4",
          4294 => x"16705381",
          4295 => x"17335259",
          4296 => x"faa23f81",
          4297 => x"dccc087a",
          4298 => x"2e098106",
          4299 => x"b73881dc",
          4300 => x"cc088317",
          4301 => x"34b01608",
          4302 => x"70a41808",
          4303 => x"319c1808",
          4304 => x"59565874",
          4305 => x"77279f38",
          4306 => x"82163355",
          4307 => x"74822e09",
          4308 => x"81069338",
          4309 => x"81547618",
          4310 => x"53785281",
          4311 => x"163351f9",
          4312 => x"e33f8339",
          4313 => x"815a7981",
          4314 => x"dccc0c8b",
          4315 => x"3d0d04fa",
          4316 => x"3d0d787a",
          4317 => x"56568057",
          4318 => x"74b01708",
          4319 => x"2eaf3875",
          4320 => x"51fefc3f",
          4321 => x"81dccc08",
          4322 => x"5781dccc",
          4323 => x"089f3881",
          4324 => x"547453b4",
          4325 => x"16528116",
          4326 => x"3351f7be",
          4327 => x"3f81dccc",
          4328 => x"08802e85",
          4329 => x"38ff5581",
          4330 => x"5774b017",
          4331 => x"0c7681dc",
          4332 => x"cc0c883d",
          4333 => x"0d04f83d",
          4334 => x"0d7a7052",
          4335 => x"57fec03f",
          4336 => x"81dccc08",
          4337 => x"5881dccc",
          4338 => x"08819138",
          4339 => x"76335574",
          4340 => x"832e0981",
          4341 => x"0680f038",
          4342 => x"84173359",
          4343 => x"78812e09",
          4344 => x"810680e3",
          4345 => x"38848053",
          4346 => x"81dccc08",
          4347 => x"52b41770",
          4348 => x"5256fd91",
          4349 => x"3f82d4d5",
          4350 => x"5284b217",
          4351 => x"51fc963f",
          4352 => x"848b85a4",
          4353 => x"d2527551",
          4354 => x"fca93f86",
          4355 => x"8a85e4f2",
          4356 => x"52849817",
          4357 => x"51fc9c3f",
          4358 => x"90170852",
          4359 => x"849c1751",
          4360 => x"fc913f8c",
          4361 => x"17085284",
          4362 => x"a01751fc",
          4363 => x"863fa017",
          4364 => x"08810570",
          4365 => x"b0190c79",
          4366 => x"55537552",
          4367 => x"81173351",
          4368 => x"f8823f77",
          4369 => x"84183480",
          4370 => x"53805281",
          4371 => x"173351f9",
          4372 => x"d73f81dc",
          4373 => x"cc08802e",
          4374 => x"83388158",
          4375 => x"7781dccc",
          4376 => x"0c8a3d0d",
          4377 => x"04fb3d0d",
          4378 => x"77fe1a98",
          4379 => x"1208fe05",
          4380 => x"55565480",
          4381 => x"56747327",
          4382 => x"8d388a14",
          4383 => x"22757129",
          4384 => x"ac160805",
          4385 => x"57537581",
          4386 => x"dccc0c87",
          4387 => x"3d0d04f9",
          4388 => x"3d0d7a7a",
          4389 => x"70085654",
          4390 => x"57817727",
          4391 => x"81df3876",
          4392 => x"98150827",
          4393 => x"81d738ff",
          4394 => x"74335458",
          4395 => x"72822e80",
          4396 => x"f5387282",
          4397 => x"24893872",
          4398 => x"812e8d38",
          4399 => x"81bf3972",
          4400 => x"832e818e",
          4401 => x"3881b639",
          4402 => x"76812a17",
          4403 => x"70892aa4",
          4404 => x"16080553",
          4405 => x"745255fd",
          4406 => x"963f81dc",
          4407 => x"cc08819f",
          4408 => x"387483ff",
          4409 => x"0614b411",
          4410 => x"33811770",
          4411 => x"892aa418",
          4412 => x"08055576",
          4413 => x"54575753",
          4414 => x"fcf53f81",
          4415 => x"dccc0880",
          4416 => x"fe387483",
          4417 => x"ff0614b4",
          4418 => x"11337088",
          4419 => x"2b780779",
          4420 => x"81067184",
          4421 => x"2a5c5258",
          4422 => x"51537280",
          4423 => x"e238759f",
          4424 => x"ff065880",
          4425 => x"da397688",
          4426 => x"2aa41508",
          4427 => x"05527351",
          4428 => x"fcbd3f81",
          4429 => x"dccc0880",
          4430 => x"c6387610",
          4431 => x"83fe0674",
          4432 => x"05b40551",
          4433 => x"f98d3f81",
          4434 => x"dccc0883",
          4435 => x"ffff0658",
          4436 => x"ae397687",
          4437 => x"2aa41508",
          4438 => x"05527351",
          4439 => x"fc913f81",
          4440 => x"dccc089b",
          4441 => x"3876822b",
          4442 => x"83fc0674",
          4443 => x"05b40551",
          4444 => x"f8f83f81",
          4445 => x"dccc08f0",
          4446 => x"0a065883",
          4447 => x"39815877",
          4448 => x"81dccc0c",
          4449 => x"893d0d04",
          4450 => x"f83d0d7a",
          4451 => x"7c7e5a58",
          4452 => x"56825981",
          4453 => x"7727829e",
          4454 => x"38769817",
          4455 => x"08278296",
          4456 => x"38753353",
          4457 => x"72792e81",
          4458 => x"9d387279",
          4459 => x"24893872",
          4460 => x"812e8d38",
          4461 => x"82803972",
          4462 => x"832e81b8",
          4463 => x"3881f739",
          4464 => x"76812a17",
          4465 => x"70892aa4",
          4466 => x"18080553",
          4467 => x"765255fb",
          4468 => x"9e3f81dc",
          4469 => x"cc085981",
          4470 => x"dccc0881",
          4471 => x"d9387483",
          4472 => x"ff0616b4",
          4473 => x"05811678",
          4474 => x"81065956",
          4475 => x"54775376",
          4476 => x"802e8f38",
          4477 => x"77842b9f",
          4478 => x"f0067433",
          4479 => x"8f067107",
          4480 => x"51537274",
          4481 => x"34810b83",
          4482 => x"17347489",
          4483 => x"2aa41708",
          4484 => x"05527551",
          4485 => x"fad93f81",
          4486 => x"dccc0859",
          4487 => x"81dccc08",
          4488 => x"81943874",
          4489 => x"83ff0616",
          4490 => x"b4057884",
          4491 => x"2a545476",
          4492 => x"8f387788",
          4493 => x"2a743381",
          4494 => x"f006718f",
          4495 => x"06075153",
          4496 => x"72743480",
          4497 => x"ec397688",
          4498 => x"2aa41708",
          4499 => x"05527551",
          4500 => x"fa9d3f81",
          4501 => x"dccc0859",
          4502 => x"81dccc08",
          4503 => x"80d83877",
          4504 => x"83ffff06",
          4505 => x"52761083",
          4506 => x"fe067605",
          4507 => x"b40551f7",
          4508 => x"a43fbe39",
          4509 => x"76872aa4",
          4510 => x"17080552",
          4511 => x"7551f9ef",
          4512 => x"3f81dccc",
          4513 => x"085981dc",
          4514 => x"cc08ab38",
          4515 => x"77f00a06",
          4516 => x"77822b83",
          4517 => x"fc067018",
          4518 => x"b4057054",
          4519 => x"515454f6",
          4520 => x"c93f81dc",
          4521 => x"cc088f0a",
          4522 => x"06740752",
          4523 => x"7251f783",
          4524 => x"3f810b83",
          4525 => x"17347881",
          4526 => x"dccc0c8a",
          4527 => x"3d0d04f8",
          4528 => x"3d0d7a7c",
          4529 => x"7e720859",
          4530 => x"56565981",
          4531 => x"7527a438",
          4532 => x"74981708",
          4533 => x"279d3873",
          4534 => x"802eaa38",
          4535 => x"ff537352",
          4536 => x"7551fda4",
          4537 => x"3f81dccc",
          4538 => x"085481dc",
          4539 => x"cc0880f2",
          4540 => x"38933982",
          4541 => x"5480eb39",
          4542 => x"815480e6",
          4543 => x"3981dccc",
          4544 => x"085480de",
          4545 => x"39745278",
          4546 => x"51fb843f",
          4547 => x"81dccc08",
          4548 => x"5881dccc",
          4549 => x"08802e80",
          4550 => x"c73881dc",
          4551 => x"cc08812e",
          4552 => x"d23881dc",
          4553 => x"cc08ff2e",
          4554 => x"cf388053",
          4555 => x"74527551",
          4556 => x"fcd63f81",
          4557 => x"dccc08c5",
          4558 => x"38981608",
          4559 => x"fe119018",
          4560 => x"08575557",
          4561 => x"74742790",
          4562 => x"38811590",
          4563 => x"170c8416",
          4564 => x"33810754",
          4565 => x"73841734",
          4566 => x"77557678",
          4567 => x"26ffa638",
          4568 => x"80547381",
          4569 => x"dccc0c8a",
          4570 => x"3d0d04f6",
          4571 => x"3d0d7c7e",
          4572 => x"7108595b",
          4573 => x"5b799538",
          4574 => x"8c170858",
          4575 => x"77802e88",
          4576 => x"38981708",
          4577 => x"7826b238",
          4578 => x"8158ae39",
          4579 => x"79527a51",
          4580 => x"f9fd3f81",
          4581 => x"557481dc",
          4582 => x"cc082782",
          4583 => x"e03881dc",
          4584 => x"cc085581",
          4585 => x"dccc08ff",
          4586 => x"2e82d238",
          4587 => x"98170881",
          4588 => x"dccc0826",
          4589 => x"82c73879",
          4590 => x"58901708",
          4591 => x"70565473",
          4592 => x"802e82b9",
          4593 => x"38777a2e",
          4594 => x"09810680",
          4595 => x"e238811a",
          4596 => x"56981708",
          4597 => x"76268338",
          4598 => x"82567552",
          4599 => x"7a51f9af",
          4600 => x"3f805981",
          4601 => x"dccc0881",
          4602 => x"2e098106",
          4603 => x"863881dc",
          4604 => x"cc085981",
          4605 => x"dccc0809",
          4606 => x"70307072",
          4607 => x"07802570",
          4608 => x"7c0781dc",
          4609 => x"cc085451",
          4610 => x"51555573",
          4611 => x"81ef3881",
          4612 => x"dccc0880",
          4613 => x"2e95388c",
          4614 => x"17085481",
          4615 => x"74279038",
          4616 => x"73981808",
          4617 => x"27893873",
          4618 => x"58853975",
          4619 => x"80db3877",
          4620 => x"56811656",
          4621 => x"98170876",
          4622 => x"26893882",
          4623 => x"56757826",
          4624 => x"81ac3875",
          4625 => x"527a51f8",
          4626 => x"c63f81dc",
          4627 => x"cc08802e",
          4628 => x"b8388059",
          4629 => x"81dccc08",
          4630 => x"812e0981",
          4631 => x"06863881",
          4632 => x"dccc0859",
          4633 => x"81dccc08",
          4634 => x"09703070",
          4635 => x"72078025",
          4636 => x"707c0751",
          4637 => x"51555573",
          4638 => x"80f83875",
          4639 => x"782e0981",
          4640 => x"06ffae38",
          4641 => x"735580f5",
          4642 => x"39ff5375",
          4643 => x"527651f9",
          4644 => x"f73f81dc",
          4645 => x"cc0881dc",
          4646 => x"cc083070",
          4647 => x"81dccc08",
          4648 => x"07802551",
          4649 => x"55557980",
          4650 => x"2e943873",
          4651 => x"802e8f38",
          4652 => x"75537952",
          4653 => x"7651f9d0",
          4654 => x"3f81dccc",
          4655 => x"085574a5",
          4656 => x"38758c18",
          4657 => x"0c981708",
          4658 => x"fe059018",
          4659 => x"08565474",
          4660 => x"74268638",
          4661 => x"ff159018",
          4662 => x"0c841733",
          4663 => x"81075473",
          4664 => x"84183497",
          4665 => x"39ff5674",
          4666 => x"812e9038",
          4667 => x"8c398055",
          4668 => x"8c3981dc",
          4669 => x"cc085585",
          4670 => x"39815675",
          4671 => x"557481dc",
          4672 => x"cc0c8c3d",
          4673 => x"0d04f83d",
          4674 => x"0d7a7052",
          4675 => x"55f3f03f",
          4676 => x"81dccc08",
          4677 => x"58815681",
          4678 => x"dccc0880",
          4679 => x"d8387b52",
          4680 => x"7451f6c1",
          4681 => x"3f81dccc",
          4682 => x"0881dccc",
          4683 => x"08b0170c",
          4684 => x"59848053",
          4685 => x"7752b415",
          4686 => x"705257f2",
          4687 => x"c83f7756",
          4688 => x"84398116",
          4689 => x"568a1522",
          4690 => x"58757827",
          4691 => x"97388154",
          4692 => x"75195376",
          4693 => x"52811533",
          4694 => x"51ede93f",
          4695 => x"81dccc08",
          4696 => x"802edf38",
          4697 => x"8a152276",
          4698 => x"32703070",
          4699 => x"7207709f",
          4700 => x"2a535156",
          4701 => x"567581dc",
          4702 => x"cc0c8a3d",
          4703 => x"0d04f83d",
          4704 => x"0d7a7c71",
          4705 => x"08585657",
          4706 => x"74f0800a",
          4707 => x"2680f138",
          4708 => x"749f0653",
          4709 => x"7280e938",
          4710 => x"7490180c",
          4711 => x"88170854",
          4712 => x"73aa3875",
          4713 => x"33538273",
          4714 => x"278838a8",
          4715 => x"16085473",
          4716 => x"9b387485",
          4717 => x"2a53820b",
          4718 => x"8817225a",
          4719 => x"58727927",
          4720 => x"80fe38a8",
          4721 => x"16089818",
          4722 => x"0c80cd39",
          4723 => x"8a162270",
          4724 => x"892b5458",
          4725 => x"727526b2",
          4726 => x"38735276",
          4727 => x"51f5b03f",
          4728 => x"81dccc08",
          4729 => x"5481dccc",
          4730 => x"08ff2ebd",
          4731 => x"38810b81",
          4732 => x"dccc0827",
          4733 => x"8b389816",
          4734 => x"0881dccc",
          4735 => x"08268538",
          4736 => x"8258bd39",
          4737 => x"74733155",
          4738 => x"cb397352",
          4739 => x"7551f4d5",
          4740 => x"3f81dccc",
          4741 => x"0898180c",
          4742 => x"7394180c",
          4743 => x"98170853",
          4744 => x"82587280",
          4745 => x"2e9a3885",
          4746 => x"39815894",
          4747 => x"3974892a",
          4748 => x"1398180c",
          4749 => x"7483ff06",
          4750 => x"16b4059c",
          4751 => x"180c8058",
          4752 => x"7781dccc",
          4753 => x"0c8a3d0d",
          4754 => x"04f83d0d",
          4755 => x"7a700890",
          4756 => x"1208a005",
          4757 => x"595754f0",
          4758 => x"800a7727",
          4759 => x"8638800b",
          4760 => x"98150c98",
          4761 => x"14085384",
          4762 => x"5572802e",
          4763 => x"81cb3876",
          4764 => x"83ff0658",
          4765 => x"7781b538",
          4766 => x"81139815",
          4767 => x"0c941408",
          4768 => x"55749238",
          4769 => x"76852a88",
          4770 => x"17225653",
          4771 => x"74732681",
          4772 => x"9b3880c0",
          4773 => x"398a1622",
          4774 => x"ff057789",
          4775 => x"2a065372",
          4776 => x"818a3874",
          4777 => x"527351f3",
          4778 => x"e63f81dc",
          4779 => x"cc085382",
          4780 => x"55810b81",
          4781 => x"dccc0827",
          4782 => x"80ff3881",
          4783 => x"5581dccc",
          4784 => x"08ff2e80",
          4785 => x"f4389816",
          4786 => x"0881dccc",
          4787 => x"082680ca",
          4788 => x"387b8a38",
          4789 => x"7798150c",
          4790 => x"845580dd",
          4791 => x"39941408",
          4792 => x"527351f9",
          4793 => x"863f81dc",
          4794 => x"cc085387",
          4795 => x"5581dccc",
          4796 => x"08802e80",
          4797 => x"c4388255",
          4798 => x"81dccc08",
          4799 => x"812eba38",
          4800 => x"815581dc",
          4801 => x"cc08ff2e",
          4802 => x"b03881dc",
          4803 => x"cc085275",
          4804 => x"51fbf33f",
          4805 => x"81dccc08",
          4806 => x"a0387294",
          4807 => x"150c7252",
          4808 => x"7551f2c1",
          4809 => x"3f81dccc",
          4810 => x"0898150c",
          4811 => x"7690150c",
          4812 => x"7716b405",
          4813 => x"9c150c80",
          4814 => x"557481dc",
          4815 => x"cc0c8a3d",
          4816 => x"0d04f73d",
          4817 => x"0d7b7d71",
          4818 => x"085b5b57",
          4819 => x"80527651",
          4820 => x"fcac3f81",
          4821 => x"dccc0854",
          4822 => x"81dccc08",
          4823 => x"80ec3881",
          4824 => x"dccc0856",
          4825 => x"98170852",
          4826 => x"7851f083",
          4827 => x"3f81dccc",
          4828 => x"085481dc",
          4829 => x"cc0880d2",
          4830 => x"3881dccc",
          4831 => x"089c1808",
          4832 => x"70335154",
          4833 => x"587281e5",
          4834 => x"2e098106",
          4835 => x"83388158",
          4836 => x"81dccc08",
          4837 => x"55728338",
          4838 => x"81557775",
          4839 => x"07537280",
          4840 => x"2e8e3881",
          4841 => x"1656757a",
          4842 => x"2e098106",
          4843 => x"8838a539",
          4844 => x"81dccc08",
          4845 => x"56815276",
          4846 => x"51fd8e3f",
          4847 => x"81dccc08",
          4848 => x"5481dccc",
          4849 => x"08802eff",
          4850 => x"9b387384",
          4851 => x"2e098106",
          4852 => x"83388754",
          4853 => x"7381dccc",
          4854 => x"0c8b3d0d",
          4855 => x"04fd3d0d",
          4856 => x"769a1152",
          4857 => x"54ebec3f",
          4858 => x"81dccc08",
          4859 => x"83ffff06",
          4860 => x"76703351",
          4861 => x"53537183",
          4862 => x"2e098106",
          4863 => x"90389414",
          4864 => x"51ebd03f",
          4865 => x"81dccc08",
          4866 => x"902b7307",
          4867 => x"537281dc",
          4868 => x"cc0c853d",
          4869 => x"0d04fc3d",
          4870 => x"0d777970",
          4871 => x"83ffff06",
          4872 => x"549a1253",
          4873 => x"5555ebed",
          4874 => x"3f767033",
          4875 => x"51537283",
          4876 => x"2e098106",
          4877 => x"8b387390",
          4878 => x"2a529415",
          4879 => x"51ebd63f",
          4880 => x"863d0d04",
          4881 => x"f73d0d7b",
          4882 => x"7d5b5584",
          4883 => x"75085a58",
          4884 => x"98150880",
          4885 => x"2e818a38",
          4886 => x"98150852",
          4887 => x"7851ee8f",
          4888 => x"3f81dccc",
          4889 => x"085881dc",
          4890 => x"cc0880f5",
          4891 => x"389c1508",
          4892 => x"70335553",
          4893 => x"73863884",
          4894 => x"5880e639",
          4895 => x"8b133370",
          4896 => x"bf067081",
          4897 => x"ff065851",
          4898 => x"53728616",
          4899 => x"3481dccc",
          4900 => x"08537381",
          4901 => x"e52e8338",
          4902 => x"815373ae",
          4903 => x"2ea93881",
          4904 => x"70740654",
          4905 => x"5772802e",
          4906 => x"9e38758f",
          4907 => x"2e993881",
          4908 => x"dccc0876",
          4909 => x"df065454",
          4910 => x"72882e09",
          4911 => x"81068338",
          4912 => x"7654737a",
          4913 => x"2ea03880",
          4914 => x"527451fa",
          4915 => x"fc3f81dc",
          4916 => x"cc085881",
          4917 => x"dccc0889",
          4918 => x"38981508",
          4919 => x"fefa3886",
          4920 => x"39800b98",
          4921 => x"160c7781",
          4922 => x"dccc0c8b",
          4923 => x"3d0d04fb",
          4924 => x"3d0d7770",
          4925 => x"08575481",
          4926 => x"527351fc",
          4927 => x"c53f81dc",
          4928 => x"cc085581",
          4929 => x"dccc08b4",
          4930 => x"38981408",
          4931 => x"527551ec",
          4932 => x"de3f81dc",
          4933 => x"cc085581",
          4934 => x"dccc08a0",
          4935 => x"38a05381",
          4936 => x"dccc0852",
          4937 => x"9c140851",
          4938 => x"eadb3f8b",
          4939 => x"53a01452",
          4940 => x"9c140851",
          4941 => x"eaac3f81",
          4942 => x"0b831734",
          4943 => x"7481dccc",
          4944 => x"0c873d0d",
          4945 => x"04fd3d0d",
          4946 => x"75700898",
          4947 => x"12085470",
          4948 => x"535553ec",
          4949 => x"9a3f81dc",
          4950 => x"cc088d38",
          4951 => x"9c130853",
          4952 => x"e5733481",
          4953 => x"0b831534",
          4954 => x"853d0d04",
          4955 => x"fa3d0d78",
          4956 => x"7a575780",
          4957 => x"0b891734",
          4958 => x"98170880",
          4959 => x"2e818238",
          4960 => x"80708918",
          4961 => x"5555559c",
          4962 => x"17081470",
          4963 => x"33811656",
          4964 => x"515271a0",
          4965 => x"2ea83871",
          4966 => x"852e0981",
          4967 => x"06843881",
          4968 => x"e5527389",
          4969 => x"2e098106",
          4970 => x"8b38ae73",
          4971 => x"70810555",
          4972 => x"34811555",
          4973 => x"71737081",
          4974 => x"05553481",
          4975 => x"15558a74",
          4976 => x"27c53875",
          4977 => x"15880552",
          4978 => x"800b8113",
          4979 => x"349c1708",
          4980 => x"528b1233",
          4981 => x"8817349c",
          4982 => x"17089c11",
          4983 => x"5252e88a",
          4984 => x"3f81dccc",
          4985 => x"08760c96",
          4986 => x"1251e7e7",
          4987 => x"3f81dccc",
          4988 => x"08861723",
          4989 => x"981251e7",
          4990 => x"da3f81dc",
          4991 => x"cc088417",
          4992 => x"23883d0d",
          4993 => x"04f33d0d",
          4994 => x"7f70085e",
          4995 => x"5b806170",
          4996 => x"33515555",
          4997 => x"73af2e83",
          4998 => x"38815573",
          4999 => x"80dc2e91",
          5000 => x"3874802e",
          5001 => x"8c38941d",
          5002 => x"08881c0c",
          5003 => x"aa398115",
          5004 => x"41806170",
          5005 => x"33565656",
          5006 => x"73af2e09",
          5007 => x"81068338",
          5008 => x"81567380",
          5009 => x"dc327030",
          5010 => x"70802578",
          5011 => x"07515154",
          5012 => x"73dc3873",
          5013 => x"881c0c60",
          5014 => x"70335154",
          5015 => x"739f2696",
          5016 => x"38ff800b",
          5017 => x"ab1c3480",
          5018 => x"527a51f6",
          5019 => x"913f81dc",
          5020 => x"cc085585",
          5021 => x"9839913d",
          5022 => x"61a01d5c",
          5023 => x"5a5e8b53",
          5024 => x"a0527951",
          5025 => x"e7ff3f80",
          5026 => x"70595788",
          5027 => x"7933555c",
          5028 => x"73ae2e09",
          5029 => x"810680d4",
          5030 => x"38781870",
          5031 => x"33811a71",
          5032 => x"ae327030",
          5033 => x"709f2a73",
          5034 => x"82260751",
          5035 => x"51535a57",
          5036 => x"54738c38",
          5037 => x"79175475",
          5038 => x"74348117",
          5039 => x"57db3975",
          5040 => x"af327030",
          5041 => x"709f2a51",
          5042 => x"51547580",
          5043 => x"dc2e8c38",
          5044 => x"73802e87",
          5045 => x"3875a026",
          5046 => x"82bd3877",
          5047 => x"197e0ca4",
          5048 => x"54a07627",
          5049 => x"82bd38a0",
          5050 => x"5482b839",
          5051 => x"78187033",
          5052 => x"811a5a57",
          5053 => x"54a07627",
          5054 => x"81fc3875",
          5055 => x"af327030",
          5056 => x"7780dc32",
          5057 => x"70307280",
          5058 => x"25718025",
          5059 => x"07515156",
          5060 => x"51557380",
          5061 => x"2eac3884",
          5062 => x"39811858",
          5063 => x"80781a70",
          5064 => x"33515555",
          5065 => x"73af2e09",
          5066 => x"81068338",
          5067 => x"81557380",
          5068 => x"dc327030",
          5069 => x"70802577",
          5070 => x"07515154",
          5071 => x"73db3881",
          5072 => x"b53975ae",
          5073 => x"2e098106",
          5074 => x"83388154",
          5075 => x"767c2774",
          5076 => x"07547380",
          5077 => x"2ea2387b",
          5078 => x"8b327030",
          5079 => x"77ae3270",
          5080 => x"30728025",
          5081 => x"719f2a07",
          5082 => x"53515651",
          5083 => x"557481a7",
          5084 => x"3888578b",
          5085 => x"5cfef539",
          5086 => x"75982b54",
          5087 => x"7380258c",
          5088 => x"387580ff",
          5089 => x"0681cc9c",
          5090 => x"11335754",
          5091 => x"7551e6e1",
          5092 => x"3f81dccc",
          5093 => x"08802eb2",
          5094 => x"38781870",
          5095 => x"33811a71",
          5096 => x"545a5654",
          5097 => x"e6d23f81",
          5098 => x"dccc0880",
          5099 => x"2e80e838",
          5100 => x"ff1c5476",
          5101 => x"742780df",
          5102 => x"38791754",
          5103 => x"75743481",
          5104 => x"177a1155",
          5105 => x"57747434",
          5106 => x"a7397552",
          5107 => x"81cbbc51",
          5108 => x"e5fe3f81",
          5109 => x"dccc08bf",
          5110 => x"38ff9f16",
          5111 => x"54739926",
          5112 => x"8938e016",
          5113 => x"7081ff06",
          5114 => x"57547917",
          5115 => x"54757434",
          5116 => x"811757fd",
          5117 => x"f7397719",
          5118 => x"7e0c7680",
          5119 => x"2e993879",
          5120 => x"33547381",
          5121 => x"e52e0981",
          5122 => x"06843885",
          5123 => x"7a348454",
          5124 => x"a076278f",
          5125 => x"388b3986",
          5126 => x"5581f239",
          5127 => x"845680f3",
          5128 => x"39805473",
          5129 => x"8b1b3480",
          5130 => x"7b085852",
          5131 => x"7a51f2ce",
          5132 => x"3f81dccc",
          5133 => x"085681dc",
          5134 => x"cc0880d7",
          5135 => x"38981b08",
          5136 => x"527651e6",
          5137 => x"aa3f81dc",
          5138 => x"cc085681",
          5139 => x"dccc0880",
          5140 => x"c2389c1b",
          5141 => x"08703355",
          5142 => x"5573802e",
          5143 => x"ffbe388b",
          5144 => x"1533bf06",
          5145 => x"5473861c",
          5146 => x"348b1533",
          5147 => x"70832a70",
          5148 => x"81065155",
          5149 => x"58739238",
          5150 => x"8b537952",
          5151 => x"7451e49f",
          5152 => x"3f81dccc",
          5153 => x"08802e8b",
          5154 => x"3875527a",
          5155 => x"51f3ba3f",
          5156 => x"ff9f3975",
          5157 => x"ab1c3357",
          5158 => x"5574802e",
          5159 => x"bb387484",
          5160 => x"2e098106",
          5161 => x"80e73875",
          5162 => x"852a7081",
          5163 => x"0677822a",
          5164 => x"58515473",
          5165 => x"802e9638",
          5166 => x"75810654",
          5167 => x"73802efb",
          5168 => x"b538ff80",
          5169 => x"0bab1c34",
          5170 => x"805580c1",
          5171 => x"39758106",
          5172 => x"5473ba38",
          5173 => x"8555b639",
          5174 => x"75822a70",
          5175 => x"81065154",
          5176 => x"73ab3886",
          5177 => x"1b337084",
          5178 => x"2a708106",
          5179 => x"51555573",
          5180 => x"802ee138",
          5181 => x"901b0883",
          5182 => x"ff061db4",
          5183 => x"05527c51",
          5184 => x"f5db3f81",
          5185 => x"dccc0888",
          5186 => x"1c0cfaea",
          5187 => x"397481dc",
          5188 => x"cc0c8f3d",
          5189 => x"0d04f63d",
          5190 => x"0d7c5bff",
          5191 => x"7b087071",
          5192 => x"7355595c",
          5193 => x"55597380",
          5194 => x"2e81c638",
          5195 => x"75708105",
          5196 => x"573370a0",
          5197 => x"26525271",
          5198 => x"ba2e8d38",
          5199 => x"70ee3871",
          5200 => x"ba2e0981",
          5201 => x"0681a538",
          5202 => x"7333d011",
          5203 => x"7081ff06",
          5204 => x"51525370",
          5205 => x"89269138",
          5206 => x"82147381",
          5207 => x"ff06d005",
          5208 => x"56527176",
          5209 => x"2e80f738",
          5210 => x"800b81cc",
          5211 => x"8c595577",
          5212 => x"087a5557",
          5213 => x"76708105",
          5214 => x"58337470",
          5215 => x"81055633",
          5216 => x"ff9f1253",
          5217 => x"53537099",
          5218 => x"268938e0",
          5219 => x"137081ff",
          5220 => x"065451ff",
          5221 => x"9f125170",
          5222 => x"99268938",
          5223 => x"e0127081",
          5224 => x"ff065351",
          5225 => x"7230709f",
          5226 => x"2a515172",
          5227 => x"722e0981",
          5228 => x"06853870",
          5229 => x"ffbe3872",
          5230 => x"30747732",
          5231 => x"70307072",
          5232 => x"079f2a73",
          5233 => x"9f2a0753",
          5234 => x"54545170",
          5235 => x"802e8f38",
          5236 => x"81158419",
          5237 => x"59558375",
          5238 => x"25ff9438",
          5239 => x"8b397483",
          5240 => x"24863874",
          5241 => x"767c0c59",
          5242 => x"78518639",
          5243 => x"81dcfc33",
          5244 => x"517081dc",
          5245 => x"cc0c8c3d",
          5246 => x"0d04fa3d",
          5247 => x"0d785680",
          5248 => x"0b831734",
          5249 => x"ff0bb017",
          5250 => x"0c795275",
          5251 => x"51e2e03f",
          5252 => x"845581dc",
          5253 => x"cc088180",
          5254 => x"3884b216",
          5255 => x"51dfb43f",
          5256 => x"81dccc08",
          5257 => x"83ffff06",
          5258 => x"54835573",
          5259 => x"82d4d52e",
          5260 => x"09810680",
          5261 => x"e338800b",
          5262 => x"b4173356",
          5263 => x"577481e9",
          5264 => x"2e098106",
          5265 => x"83388157",
          5266 => x"7481eb32",
          5267 => x"70307080",
          5268 => x"25790751",
          5269 => x"5154738a",
          5270 => x"387481e8",
          5271 => x"2e098106",
          5272 => x"b5388353",
          5273 => x"81cbcc52",
          5274 => x"80ea1651",
          5275 => x"e0b13f81",
          5276 => x"dccc0855",
          5277 => x"81dccc08",
          5278 => x"802e9d38",
          5279 => x"855381cb",
          5280 => x"d0528186",
          5281 => x"1651e097",
          5282 => x"3f81dccc",
          5283 => x"085581dc",
          5284 => x"cc08802e",
          5285 => x"83388255",
          5286 => x"7481dccc",
          5287 => x"0c883d0d",
          5288 => x"04f23d0d",
          5289 => x"61028405",
          5290 => x"80cb0533",
          5291 => x"58558075",
          5292 => x"0c6051fc",
          5293 => x"e13f81dc",
          5294 => x"cc08588b",
          5295 => x"56800b81",
          5296 => x"dccc0824",
          5297 => x"86fc3881",
          5298 => x"dccc0884",
          5299 => x"2981dce8",
          5300 => x"05700855",
          5301 => x"538c5673",
          5302 => x"802e86e6",
          5303 => x"3873750c",
          5304 => x"7681fe06",
          5305 => x"74335457",
          5306 => x"72802eae",
          5307 => x"38811433",
          5308 => x"51d7ca3f",
          5309 => x"81dccc08",
          5310 => x"81ff0670",
          5311 => x"81065455",
          5312 => x"72983876",
          5313 => x"802e86b8",
          5314 => x"3874822a",
          5315 => x"70810651",
          5316 => x"538a5672",
          5317 => x"86ac3886",
          5318 => x"a7398074",
          5319 => x"34778115",
          5320 => x"34815281",
          5321 => x"143351d7",
          5322 => x"b23f81dc",
          5323 => x"cc0881ff",
          5324 => x"06708106",
          5325 => x"54558356",
          5326 => x"72868738",
          5327 => x"76802e8f",
          5328 => x"3874822a",
          5329 => x"70810651",
          5330 => x"538a5672",
          5331 => x"85f43880",
          5332 => x"70537452",
          5333 => x"5bfda33f",
          5334 => x"81dccc08",
          5335 => x"81ff0657",
          5336 => x"76822e09",
          5337 => x"810680e2",
          5338 => x"388c3d74",
          5339 => x"56588356",
          5340 => x"83f61533",
          5341 => x"70585372",
          5342 => x"802e8d38",
          5343 => x"83fa1551",
          5344 => x"dce83f81",
          5345 => x"dccc0857",
          5346 => x"76787084",
          5347 => x"055a0cff",
          5348 => x"16901656",
          5349 => x"56758025",
          5350 => x"d738800b",
          5351 => x"8d3d5456",
          5352 => x"72708405",
          5353 => x"54085b83",
          5354 => x"577a802e",
          5355 => x"95387a52",
          5356 => x"7351fcc6",
          5357 => x"3f81dccc",
          5358 => x"0881ff06",
          5359 => x"57817727",
          5360 => x"89388116",
          5361 => x"56837627",
          5362 => x"d7388156",
          5363 => x"76842e84",
          5364 => x"f1388d56",
          5365 => x"76812684",
          5366 => x"e938bf14",
          5367 => x"51dbf43f",
          5368 => x"81dccc08",
          5369 => x"83ffff06",
          5370 => x"53728480",
          5371 => x"2e098106",
          5372 => x"84d03880",
          5373 => x"ca1451db",
          5374 => x"da3f81dc",
          5375 => x"cc0883ff",
          5376 => x"ff065877",
          5377 => x"8d3880d8",
          5378 => x"1451dbde",
          5379 => x"3f81dccc",
          5380 => x"0858779c",
          5381 => x"150c80c4",
          5382 => x"14338215",
          5383 => x"3480c414",
          5384 => x"33ff1170",
          5385 => x"81ff0651",
          5386 => x"54558d56",
          5387 => x"72812684",
          5388 => x"91387481",
          5389 => x"ff067871",
          5390 => x"2980c116",
          5391 => x"33525953",
          5392 => x"728a1523",
          5393 => x"72802e8b",
          5394 => x"38ff1373",
          5395 => x"06537280",
          5396 => x"2e86388d",
          5397 => x"5683eb39",
          5398 => x"80c51451",
          5399 => x"daf53f81",
          5400 => x"dccc0853",
          5401 => x"81dccc08",
          5402 => x"88152372",
          5403 => x"8f06578d",
          5404 => x"567683ce",
          5405 => x"3880c714",
          5406 => x"51dad83f",
          5407 => x"81dccc08",
          5408 => x"83ffff06",
          5409 => x"55748d38",
          5410 => x"80d41451",
          5411 => x"dadc3f81",
          5412 => x"dccc0855",
          5413 => x"80c21451",
          5414 => x"dab93f81",
          5415 => x"dccc0883",
          5416 => x"ffff0653",
          5417 => x"8d567280",
          5418 => x"2e839738",
          5419 => x"88142278",
          5420 => x"1471842a",
          5421 => x"055a5a78",
          5422 => x"75268386",
          5423 => x"388a1422",
          5424 => x"52747931",
          5425 => x"51ffadb1",
          5426 => x"3f81dccc",
          5427 => x"085581dc",
          5428 => x"cc08802e",
          5429 => x"82ec3881",
          5430 => x"dccc0880",
          5431 => x"fffffff5",
          5432 => x"26833883",
          5433 => x"577483ff",
          5434 => x"f5268338",
          5435 => x"8257749f",
          5436 => x"f5268538",
          5437 => x"81578939",
          5438 => x"8d567680",
          5439 => x"2e82c338",
          5440 => x"82157098",
          5441 => x"160c7ba0",
          5442 => x"160c731c",
          5443 => x"70a4170c",
          5444 => x"7a1dac17",
          5445 => x"0c545576",
          5446 => x"832e0981",
          5447 => x"06af3880",
          5448 => x"de1451d9",
          5449 => x"ae3f81dc",
          5450 => x"cc0883ff",
          5451 => x"ff06538d",
          5452 => x"5672828e",
          5453 => x"3879828a",
          5454 => x"3880e014",
          5455 => x"51d9ab3f",
          5456 => x"81dccc08",
          5457 => x"a8150c74",
          5458 => x"822b53a2",
          5459 => x"398d5679",
          5460 => x"802e81ee",
          5461 => x"387713a8",
          5462 => x"150c7415",
          5463 => x"5376822e",
          5464 => x"8d387410",
          5465 => x"1570812a",
          5466 => x"76810605",
          5467 => x"515383ff",
          5468 => x"13892a53",
          5469 => x"8d56729c",
          5470 => x"15082681",
          5471 => x"c538ff0b",
          5472 => x"90150cff",
          5473 => x"0b8c150c",
          5474 => x"ff800b84",
          5475 => x"15347683",
          5476 => x"2e098106",
          5477 => x"81923880",
          5478 => x"e41451d8",
          5479 => x"b63f81dc",
          5480 => x"cc0883ff",
          5481 => x"ff065372",
          5482 => x"812e0981",
          5483 => x"0680f938",
          5484 => x"811b5273",
          5485 => x"51dbb83f",
          5486 => x"81dccc08",
          5487 => x"80ea3881",
          5488 => x"dccc0884",
          5489 => x"153484b2",
          5490 => x"1451d887",
          5491 => x"3f81dccc",
          5492 => x"0883ffff",
          5493 => x"06537282",
          5494 => x"d4d52e09",
          5495 => x"810680c8",
          5496 => x"38b41451",
          5497 => x"d8843f81",
          5498 => x"dccc0884",
          5499 => x"8b85a4d2",
          5500 => x"2e098106",
          5501 => x"b3388498",
          5502 => x"1451d7ee",
          5503 => x"3f81dccc",
          5504 => x"08868a85",
          5505 => x"e4f22e09",
          5506 => x"81069d38",
          5507 => x"849c1451",
          5508 => x"d7d83f81",
          5509 => x"dccc0890",
          5510 => x"150c84a0",
          5511 => x"1451d7ca",
          5512 => x"3f81dccc",
          5513 => x"088c150c",
          5514 => x"76743481",
          5515 => x"dcf82281",
          5516 => x"05537281",
          5517 => x"dcf82372",
          5518 => x"86152380",
          5519 => x"0b94150c",
          5520 => x"80567581",
          5521 => x"dccc0c90",
          5522 => x"3d0d04fb",
          5523 => x"3d0d7754",
          5524 => x"89557380",
          5525 => x"2eb93873",
          5526 => x"08537280",
          5527 => x"2eb13872",
          5528 => x"33527180",
          5529 => x"2ea93886",
          5530 => x"13228415",
          5531 => x"22575271",
          5532 => x"762e0981",
          5533 => x"06993881",
          5534 => x"133351d0",
          5535 => x"c03f81dc",
          5536 => x"cc088106",
          5537 => x"52718838",
          5538 => x"71740854",
          5539 => x"55833980",
          5540 => x"53787371",
          5541 => x"0c527481",
          5542 => x"dccc0c87",
          5543 => x"3d0d04fa",
          5544 => x"3d0d02ab",
          5545 => x"05337a58",
          5546 => x"893dfc05",
          5547 => x"5256f4e6",
          5548 => x"3f8b5480",
          5549 => x"0b81dccc",
          5550 => x"0824bc38",
          5551 => x"81dccc08",
          5552 => x"842981dc",
          5553 => x"e8057008",
          5554 => x"55557380",
          5555 => x"2e843880",
          5556 => x"74347854",
          5557 => x"73802e84",
          5558 => x"38807434",
          5559 => x"78750c75",
          5560 => x"5475802e",
          5561 => x"92388053",
          5562 => x"893d7053",
          5563 => x"840551f7",
          5564 => x"b03f81dc",
          5565 => x"cc085473",
          5566 => x"81dccc0c",
          5567 => x"883d0d04",
          5568 => x"eb3d0d67",
          5569 => x"02840580",
          5570 => x"e7053359",
          5571 => x"59895478",
          5572 => x"802e84c8",
          5573 => x"3877bf06",
          5574 => x"7054983d",
          5575 => x"d0055399",
          5576 => x"3d840552",
          5577 => x"58f6fa3f",
          5578 => x"81dccc08",
          5579 => x"5581dccc",
          5580 => x"0884a438",
          5581 => x"7a5c6852",
          5582 => x"8c3d7052",
          5583 => x"56edc63f",
          5584 => x"81dccc08",
          5585 => x"5581dccc",
          5586 => x"08923802",
          5587 => x"80d70533",
          5588 => x"70982b55",
          5589 => x"57738025",
          5590 => x"83388655",
          5591 => x"779c0654",
          5592 => x"73802e81",
          5593 => x"ab387480",
          5594 => x"2e953874",
          5595 => x"842e0981",
          5596 => x"06aa3875",
          5597 => x"51eaf83f",
          5598 => x"81dccc08",
          5599 => x"559e3902",
          5600 => x"b2053391",
          5601 => x"06547381",
          5602 => x"b8387782",
          5603 => x"2a708106",
          5604 => x"51547380",
          5605 => x"2e8e3888",
          5606 => x"5583bc39",
          5607 => x"77880758",
          5608 => x"7483b438",
          5609 => x"77832a70",
          5610 => x"81065154",
          5611 => x"73802e81",
          5612 => x"af386252",
          5613 => x"7a51e8a5",
          5614 => x"3f81dccc",
          5615 => x"08568288",
          5616 => x"b20a5262",
          5617 => x"8e0551d4",
          5618 => x"ea3f6254",
          5619 => x"a00b8b15",
          5620 => x"34805362",
          5621 => x"527a51e8",
          5622 => x"bd3f8052",
          5623 => x"629c0551",
          5624 => x"d4d13f7a",
          5625 => x"54810b83",
          5626 => x"15347580",
          5627 => x"2e80f138",
          5628 => x"7ab01108",
          5629 => x"51548053",
          5630 => x"7552973d",
          5631 => x"d40551dd",
          5632 => x"be3f81dc",
          5633 => x"cc085581",
          5634 => x"dccc0882",
          5635 => x"ca38b739",
          5636 => x"7482c438",
          5637 => x"02b20533",
          5638 => x"70842a70",
          5639 => x"81065155",
          5640 => x"5673802e",
          5641 => x"86388455",
          5642 => x"82ad3977",
          5643 => x"812a7081",
          5644 => x"06515473",
          5645 => x"802ea938",
          5646 => x"75810654",
          5647 => x"73802ea0",
          5648 => x"38875582",
          5649 => x"92397352",
          5650 => x"7a51d6a3",
          5651 => x"3f81dccc",
          5652 => x"087bff18",
          5653 => x"8c120c55",
          5654 => x"5581dccc",
          5655 => x"0881f838",
          5656 => x"77832a70",
          5657 => x"81065154",
          5658 => x"73802e86",
          5659 => x"387780c0",
          5660 => x"07587ab0",
          5661 => x"1108a01b",
          5662 => x"0c63a41b",
          5663 => x"0c635370",
          5664 => x"5257e6d9",
          5665 => x"3f81dccc",
          5666 => x"0881dccc",
          5667 => x"08881b0c",
          5668 => x"639c0552",
          5669 => x"5ad2d33f",
          5670 => x"81dccc08",
          5671 => x"81dccc08",
          5672 => x"8c1b0c77",
          5673 => x"7a0c5686",
          5674 => x"1722841a",
          5675 => x"2377901a",
          5676 => x"34800b91",
          5677 => x"1a34800b",
          5678 => x"9c1a0c80",
          5679 => x"0b941a0c",
          5680 => x"77852a70",
          5681 => x"81065154",
          5682 => x"73802e81",
          5683 => x"8d3881dc",
          5684 => x"cc08802e",
          5685 => x"81843881",
          5686 => x"dccc0894",
          5687 => x"1a0c8a17",
          5688 => x"2270892b",
          5689 => x"7b525957",
          5690 => x"a8397652",
          5691 => x"7851d79f",
          5692 => x"3f81dccc",
          5693 => x"085781dc",
          5694 => x"cc088126",
          5695 => x"83388255",
          5696 => x"81dccc08",
          5697 => x"ff2e0981",
          5698 => x"06833879",
          5699 => x"55757831",
          5700 => x"56743070",
          5701 => x"76078025",
          5702 => x"51547776",
          5703 => x"278a3881",
          5704 => x"70750655",
          5705 => x"5a73c338",
          5706 => x"76981a0c",
          5707 => x"74a93875",
          5708 => x"83ff0654",
          5709 => x"73802ea2",
          5710 => x"3876527a",
          5711 => x"51d6a63f",
          5712 => x"81dccc08",
          5713 => x"85388255",
          5714 => x"8e397589",
          5715 => x"2a81dccc",
          5716 => x"08059c1a",
          5717 => x"0c843980",
          5718 => x"790c7454",
          5719 => x"7381dccc",
          5720 => x"0c973d0d",
          5721 => x"04f23d0d",
          5722 => x"60636564",
          5723 => x"40405d59",
          5724 => x"807e0c90",
          5725 => x"3dfc0552",
          5726 => x"7851f9cf",
          5727 => x"3f81dccc",
          5728 => x"085581dc",
          5729 => x"cc088a38",
          5730 => x"91193355",
          5731 => x"74802e86",
          5732 => x"38745682",
          5733 => x"c4399019",
          5734 => x"33810655",
          5735 => x"87567480",
          5736 => x"2e82b638",
          5737 => x"9539820b",
          5738 => x"911a3482",
          5739 => x"5682aa39",
          5740 => x"810b911a",
          5741 => x"34815682",
          5742 => x"a0398c19",
          5743 => x"08941a08",
          5744 => x"3155747c",
          5745 => x"27833874",
          5746 => x"5c7b802e",
          5747 => x"82893894",
          5748 => x"19087083",
          5749 => x"ff065656",
          5750 => x"7481b238",
          5751 => x"7e8a1122",
          5752 => x"ff057789",
          5753 => x"2a065b55",
          5754 => x"79a83875",
          5755 => x"87388819",
          5756 => x"08558f39",
          5757 => x"98190852",
          5758 => x"7851d593",
          5759 => x"3f81dccc",
          5760 => x"08558175",
          5761 => x"27ff9f38",
          5762 => x"74ff2eff",
          5763 => x"a3387498",
          5764 => x"1a0c9819",
          5765 => x"08527e51",
          5766 => x"d4cb3f81",
          5767 => x"dccc0880",
          5768 => x"2eff8338",
          5769 => x"81dccc08",
          5770 => x"1a7c892a",
          5771 => x"59577780",
          5772 => x"2e80d638",
          5773 => x"771a7f8a",
          5774 => x"1122585c",
          5775 => x"55757527",
          5776 => x"8538757a",
          5777 => x"31587754",
          5778 => x"76537c52",
          5779 => x"811b3351",
          5780 => x"ca883f81",
          5781 => x"dccc08fe",
          5782 => x"d7387e83",
          5783 => x"11335656",
          5784 => x"74802e9f",
          5785 => x"38b01608",
          5786 => x"77315574",
          5787 => x"78279438",
          5788 => x"848053b4",
          5789 => x"1652b016",
          5790 => x"08773189",
          5791 => x"2b7d0551",
          5792 => x"cfe03f77",
          5793 => x"892b56b9",
          5794 => x"39769c1a",
          5795 => x"0c941908",
          5796 => x"83ff0684",
          5797 => x"80713157",
          5798 => x"557b7627",
          5799 => x"83387b56",
          5800 => x"9c190852",
          5801 => x"7e51d1c7",
          5802 => x"3f81dccc",
          5803 => x"08fe8138",
          5804 => x"75539419",
          5805 => x"0883ff06",
          5806 => x"1fb40552",
          5807 => x"7c51cfa2",
          5808 => x"3f7b7631",
          5809 => x"7e08177f",
          5810 => x"0c761e94",
          5811 => x"1b081894",
          5812 => x"1c0c5e5c",
          5813 => x"fdf33980",
          5814 => x"567581dc",
          5815 => x"cc0c903d",
          5816 => x"0d04f23d",
          5817 => x"0d606365",
          5818 => x"6440405d",
          5819 => x"58807e0c",
          5820 => x"903dfc05",
          5821 => x"527751f6",
          5822 => x"d23f81dc",
          5823 => x"cc085581",
          5824 => x"dccc088a",
          5825 => x"38911833",
          5826 => x"5574802e",
          5827 => x"86387456",
          5828 => x"83b83990",
          5829 => x"18337081",
          5830 => x"2a708106",
          5831 => x"51565687",
          5832 => x"5674802e",
          5833 => x"83a43895",
          5834 => x"39820b91",
          5835 => x"19348256",
          5836 => x"83983981",
          5837 => x"0b911934",
          5838 => x"8156838e",
          5839 => x"39941808",
          5840 => x"7c115656",
          5841 => x"74762784",
          5842 => x"3875095c",
          5843 => x"7b802e82",
          5844 => x"ec389418",
          5845 => x"087083ff",
          5846 => x"06565674",
          5847 => x"81fd387e",
          5848 => x"8a1122ff",
          5849 => x"0577892a",
          5850 => x"065c557a",
          5851 => x"bf38758c",
          5852 => x"38881808",
          5853 => x"55749c38",
          5854 => x"7a528539",
          5855 => x"98180852",
          5856 => x"7751d7e7",
          5857 => x"3f81dccc",
          5858 => x"085581dc",
          5859 => x"cc08802e",
          5860 => x"82ab3874",
          5861 => x"812eff91",
          5862 => x"3874ff2e",
          5863 => x"ff953874",
          5864 => x"98190c88",
          5865 => x"18088538",
          5866 => x"7488190c",
          5867 => x"7e55b015",
          5868 => x"089c1908",
          5869 => x"2e098106",
          5870 => x"8d387451",
          5871 => x"cec13f81",
          5872 => x"dccc08fe",
          5873 => x"ee389818",
          5874 => x"08527e51",
          5875 => x"d1973f81",
          5876 => x"dccc0880",
          5877 => x"2efed238",
          5878 => x"81dccc08",
          5879 => x"1b7c892a",
          5880 => x"5a577880",
          5881 => x"2e80d538",
          5882 => x"781b7f8a",
          5883 => x"1122585b",
          5884 => x"55757527",
          5885 => x"8538757b",
          5886 => x"31597854",
          5887 => x"76537c52",
          5888 => x"811a3351",
          5889 => x"c8be3f81",
          5890 => x"dccc08fe",
          5891 => x"a6387eb0",
          5892 => x"11087831",
          5893 => x"56567479",
          5894 => x"279b3884",
          5895 => x"8053b016",
          5896 => x"08773189",
          5897 => x"2b7d0552",
          5898 => x"b41651cc",
          5899 => x"b53f7e55",
          5900 => x"800b8316",
          5901 => x"3478892b",
          5902 => x"5680db39",
          5903 => x"8c180894",
          5904 => x"19082693",
          5905 => x"387e51cd",
          5906 => x"b63f81dc",
          5907 => x"cc08fde3",
          5908 => x"387e77b0",
          5909 => x"120c5576",
          5910 => x"9c190c94",
          5911 => x"180883ff",
          5912 => x"06848071",
          5913 => x"3157557b",
          5914 => x"76278338",
          5915 => x"7b569c18",
          5916 => x"08527e51",
          5917 => x"cdf93f81",
          5918 => x"dccc08fd",
          5919 => x"b6387553",
          5920 => x"7c529418",
          5921 => x"0883ff06",
          5922 => x"1fb40551",
          5923 => x"cbd43f7e",
          5924 => x"55810b83",
          5925 => x"16347b76",
          5926 => x"317e0817",
          5927 => x"7f0c761e",
          5928 => x"941a0818",
          5929 => x"70941c0c",
          5930 => x"8c1b0858",
          5931 => x"585e5c74",
          5932 => x"76278338",
          5933 => x"7555748c",
          5934 => x"190cfd90",
          5935 => x"39901833",
          5936 => x"80c00755",
          5937 => x"74901934",
          5938 => x"80567581",
          5939 => x"dccc0c90",
          5940 => x"3d0d04f8",
          5941 => x"3d0d7a8b",
          5942 => x"3dfc0553",
          5943 => x"705256f2",
          5944 => x"ea3f81dc",
          5945 => x"cc085781",
          5946 => x"dccc0880",
          5947 => x"fb389016",
          5948 => x"3370862a",
          5949 => x"70810651",
          5950 => x"55557380",
          5951 => x"2e80e938",
          5952 => x"a0160852",
          5953 => x"7851cce7",
          5954 => x"3f81dccc",
          5955 => x"085781dc",
          5956 => x"cc0880d4",
          5957 => x"38a41608",
          5958 => x"8b1133a0",
          5959 => x"07555573",
          5960 => x"8b163488",
          5961 => x"16085374",
          5962 => x"52750851",
          5963 => x"dde83f8c",
          5964 => x"1608529c",
          5965 => x"1551c9fb",
          5966 => x"3f8288b2",
          5967 => x"0a529615",
          5968 => x"51c9f03f",
          5969 => x"76529215",
          5970 => x"51c9ca3f",
          5971 => x"7854810b",
          5972 => x"83153478",
          5973 => x"51ccdf3f",
          5974 => x"81dccc08",
          5975 => x"90173381",
          5976 => x"bf065557",
          5977 => x"73901734",
          5978 => x"7681dccc",
          5979 => x"0c8a3d0d",
          5980 => x"04fc3d0d",
          5981 => x"76705254",
          5982 => x"fed93f81",
          5983 => x"dccc0853",
          5984 => x"81dccc08",
          5985 => x"9c38863d",
          5986 => x"fc055273",
          5987 => x"51f1bc3f",
          5988 => x"81dccc08",
          5989 => x"5381dccc",
          5990 => x"08873881",
          5991 => x"dccc0874",
          5992 => x"0c7281dc",
          5993 => x"cc0c863d",
          5994 => x"0d04ff3d",
          5995 => x"0d843d51",
          5996 => x"e6e43f8b",
          5997 => x"52800b81",
          5998 => x"dccc0824",
          5999 => x"8b3881dc",
          6000 => x"cc0881dc",
          6001 => x"fc348052",
          6002 => x"7181dccc",
          6003 => x"0c833d0d",
          6004 => x"04ef3d0d",
          6005 => x"8053933d",
          6006 => x"d0055294",
          6007 => x"3d51e9c1",
          6008 => x"3f81dccc",
          6009 => x"085581dc",
          6010 => x"cc0880e0",
          6011 => x"38765863",
          6012 => x"52933dd4",
          6013 => x"0551e08d",
          6014 => x"3f81dccc",
          6015 => x"085581dc",
          6016 => x"cc08bc38",
          6017 => x"0280c705",
          6018 => x"3370982b",
          6019 => x"55567380",
          6020 => x"25893876",
          6021 => x"7a94120c",
          6022 => x"54b23902",
          6023 => x"a2053370",
          6024 => x"842a7081",
          6025 => x"06515556",
          6026 => x"73802e9e",
          6027 => x"38767f53",
          6028 => x"705254db",
          6029 => x"a83f81dc",
          6030 => x"cc089415",
          6031 => x"0c8e3981",
          6032 => x"dccc0884",
          6033 => x"2e098106",
          6034 => x"83388555",
          6035 => x"7481dccc",
          6036 => x"0c933d0d",
          6037 => x"04e43d0d",
          6038 => x"6f6f5b5b",
          6039 => x"807a3480",
          6040 => x"539e3dff",
          6041 => x"b805529f",
          6042 => x"3d51e8b5",
          6043 => x"3f81dccc",
          6044 => x"085781dc",
          6045 => x"cc0882fc",
          6046 => x"387b437a",
          6047 => x"7c941108",
          6048 => x"47555864",
          6049 => x"5473802e",
          6050 => x"81ed38a0",
          6051 => x"52933d70",
          6052 => x"5255d5ea",
          6053 => x"3f81dccc",
          6054 => x"085781dc",
          6055 => x"cc0882d4",
          6056 => x"3868527b",
          6057 => x"51c9c83f",
          6058 => x"81dccc08",
          6059 => x"5781dccc",
          6060 => x"0882c138",
          6061 => x"69527b51",
          6062 => x"daa33f81",
          6063 => x"dccc0845",
          6064 => x"76527451",
          6065 => x"d5b83f81",
          6066 => x"dccc0857",
          6067 => x"81dccc08",
          6068 => x"82a23880",
          6069 => x"527451da",
          6070 => x"eb3f81dc",
          6071 => x"cc085781",
          6072 => x"dccc08a4",
          6073 => x"3869527b",
          6074 => x"51d9f23f",
          6075 => x"7381dccc",
          6076 => x"082ea638",
          6077 => x"76527451",
          6078 => x"d6cf3f81",
          6079 => x"dccc0857",
          6080 => x"81dccc08",
          6081 => x"802ecc38",
          6082 => x"76842e09",
          6083 => x"81068638",
          6084 => x"825781e0",
          6085 => x"397681dc",
          6086 => x"389e3dff",
          6087 => x"bc055274",
          6088 => x"51dcc93f",
          6089 => x"76903d78",
          6090 => x"11811133",
          6091 => x"51565a56",
          6092 => x"73802e91",
          6093 => x"3802b905",
          6094 => x"55811681",
          6095 => x"16703356",
          6096 => x"565673f5",
          6097 => x"38811654",
          6098 => x"73782681",
          6099 => x"90387580",
          6100 => x"2e993878",
          6101 => x"16810555",
          6102 => x"ff186f11",
          6103 => x"ff18ff18",
          6104 => x"58585558",
          6105 => x"74337434",
          6106 => x"75ee38ff",
          6107 => x"186f1155",
          6108 => x"58af7434",
          6109 => x"fe8d3977",
          6110 => x"7b2e0981",
          6111 => x"068a38ff",
          6112 => x"186f1155",
          6113 => x"58af7434",
          6114 => x"800b81dc",
          6115 => x"fc337084",
          6116 => x"2981cc8c",
          6117 => x"05700870",
          6118 => x"33525c56",
          6119 => x"56567376",
          6120 => x"2e8d3881",
          6121 => x"16701a70",
          6122 => x"33515556",
          6123 => x"73f53882",
          6124 => x"16547378",
          6125 => x"26a73880",
          6126 => x"55747627",
          6127 => x"91387419",
          6128 => x"5473337a",
          6129 => x"7081055c",
          6130 => x"34811555",
          6131 => x"ec39ba7a",
          6132 => x"7081055c",
          6133 => x"3474ff2e",
          6134 => x"09810685",
          6135 => x"38915794",
          6136 => x"396e1881",
          6137 => x"19595473",
          6138 => x"337a7081",
          6139 => x"055c347a",
          6140 => x"7826ee38",
          6141 => x"807a3476",
          6142 => x"81dccc0c",
          6143 => x"9e3d0d04",
          6144 => x"f73d0d7b",
          6145 => x"7d8d3dfc",
          6146 => x"05547153",
          6147 => x"5755ecbb",
          6148 => x"3f81dccc",
          6149 => x"085381dc",
          6150 => x"cc0882fa",
          6151 => x"38911533",
          6152 => x"537282f2",
          6153 => x"388c1508",
          6154 => x"54737627",
          6155 => x"92389015",
          6156 => x"3370812a",
          6157 => x"70810651",
          6158 => x"54577283",
          6159 => x"38735694",
          6160 => x"15085480",
          6161 => x"7094170c",
          6162 => x"5875782e",
          6163 => x"82973879",
          6164 => x"8a112270",
          6165 => x"892b5951",
          6166 => x"5373782e",
          6167 => x"b7387652",
          6168 => x"ff1651ff",
          6169 => x"96933f81",
          6170 => x"dccc08ff",
          6171 => x"15785470",
          6172 => x"535553ff",
          6173 => x"96833f81",
          6174 => x"dccc0873",
          6175 => x"26963876",
          6176 => x"30707506",
          6177 => x"7094180c",
          6178 => x"77713198",
          6179 => x"18085758",
          6180 => x"5153b139",
          6181 => x"88150854",
          6182 => x"73a63873",
          6183 => x"527451cd",
          6184 => x"ca3f81dc",
          6185 => x"cc085481",
          6186 => x"dccc0881",
          6187 => x"2e819a38",
          6188 => x"81dccc08",
          6189 => x"ff2e819b",
          6190 => x"3881dccc",
          6191 => x"0888160c",
          6192 => x"7398160c",
          6193 => x"73802e81",
          6194 => x"9c387676",
          6195 => x"2780dc38",
          6196 => x"75773194",
          6197 => x"16081894",
          6198 => x"170c9016",
          6199 => x"3370812a",
          6200 => x"70810651",
          6201 => x"555a5672",
          6202 => x"802e9a38",
          6203 => x"73527451",
          6204 => x"ccf93f81",
          6205 => x"dccc0854",
          6206 => x"81dccc08",
          6207 => x"943881dc",
          6208 => x"cc0856a7",
          6209 => x"39735274",
          6210 => x"51c7843f",
          6211 => x"81dccc08",
          6212 => x"5473ff2e",
          6213 => x"be388174",
          6214 => x"27af3879",
          6215 => x"53739814",
          6216 => x"0827a638",
          6217 => x"7398160c",
          6218 => x"ffa03994",
          6219 => x"15081694",
          6220 => x"160c7583",
          6221 => x"ff065372",
          6222 => x"802eaa38",
          6223 => x"73527951",
          6224 => x"c6a33f81",
          6225 => x"dccc0894",
          6226 => x"38820b91",
          6227 => x"16348253",
          6228 => x"80c43981",
          6229 => x"0b911634",
          6230 => x"8153bb39",
          6231 => x"75892a81",
          6232 => x"dccc0805",
          6233 => x"58941508",
          6234 => x"548c1508",
          6235 => x"74279038",
          6236 => x"738c160c",
          6237 => x"90153380",
          6238 => x"c0075372",
          6239 => x"90163473",
          6240 => x"83ff0653",
          6241 => x"72802e8c",
          6242 => x"38779c16",
          6243 => x"082e8538",
          6244 => x"779c160c",
          6245 => x"80537281",
          6246 => x"dccc0c8b",
          6247 => x"3d0d04f9",
          6248 => x"3d0d7956",
          6249 => x"89547580",
          6250 => x"2e818a38",
          6251 => x"8053893d",
          6252 => x"fc05528a",
          6253 => x"3d840551",
          6254 => x"e1e73f81",
          6255 => x"dccc0855",
          6256 => x"81dccc08",
          6257 => x"80ea3877",
          6258 => x"760c7a52",
          6259 => x"7551d8b5",
          6260 => x"3f81dccc",
          6261 => x"085581dc",
          6262 => x"cc0880c3",
          6263 => x"38ab1633",
          6264 => x"70982b55",
          6265 => x"57807424",
          6266 => x"a2388616",
          6267 => x"3370842a",
          6268 => x"70810651",
          6269 => x"55577380",
          6270 => x"2ead389c",
          6271 => x"16085277",
          6272 => x"51d3da3f",
          6273 => x"81dccc08",
          6274 => x"88170c77",
          6275 => x"54861422",
          6276 => x"84172374",
          6277 => x"527551ce",
          6278 => x"e53f81dc",
          6279 => x"cc085574",
          6280 => x"842e0981",
          6281 => x"06853885",
          6282 => x"55863974",
          6283 => x"802e8438",
          6284 => x"80760c74",
          6285 => x"547381dc",
          6286 => x"cc0c893d",
          6287 => x"0d04fc3d",
          6288 => x"0d76873d",
          6289 => x"fc055370",
          6290 => x"5253e7ff",
          6291 => x"3f81dccc",
          6292 => x"08873881",
          6293 => x"dccc0873",
          6294 => x"0c863d0d",
          6295 => x"04fb3d0d",
          6296 => x"7779893d",
          6297 => x"fc055471",
          6298 => x"535654e7",
          6299 => x"de3f81dc",
          6300 => x"cc085381",
          6301 => x"dccc0880",
          6302 => x"df387493",
          6303 => x"3881dccc",
          6304 => x"08527351",
          6305 => x"cdf83f81",
          6306 => x"dccc0853",
          6307 => x"80ca3981",
          6308 => x"dccc0852",
          6309 => x"7351d3ac",
          6310 => x"3f81dccc",
          6311 => x"085381dc",
          6312 => x"cc08842e",
          6313 => x"09810685",
          6314 => x"38805387",
          6315 => x"3981dccc",
          6316 => x"08a63874",
          6317 => x"527351d5",
          6318 => x"b33f7252",
          6319 => x"7351cf89",
          6320 => x"3f81dccc",
          6321 => x"08843270",
          6322 => x"30707207",
          6323 => x"9f2c7081",
          6324 => x"dccc0806",
          6325 => x"51515454",
          6326 => x"7281dccc",
          6327 => x"0c873d0d",
          6328 => x"04ee3d0d",
          6329 => x"65578053",
          6330 => x"893d7053",
          6331 => x"963d5256",
          6332 => x"dfaf3f81",
          6333 => x"dccc0855",
          6334 => x"81dccc08",
          6335 => x"b2386452",
          6336 => x"7551d681",
          6337 => x"3f81dccc",
          6338 => x"085581dc",
          6339 => x"cc08a038",
          6340 => x"0280cb05",
          6341 => x"3370982b",
          6342 => x"55587380",
          6343 => x"25853886",
          6344 => x"558d3976",
          6345 => x"802e8838",
          6346 => x"76527551",
          6347 => x"d4be3f74",
          6348 => x"81dccc0c",
          6349 => x"943d0d04",
          6350 => x"f03d0d63",
          6351 => x"65555c80",
          6352 => x"53923dec",
          6353 => x"0552933d",
          6354 => x"51ded63f",
          6355 => x"81dccc08",
          6356 => x"5b81dccc",
          6357 => x"08828038",
          6358 => x"7c740c73",
          6359 => x"08981108",
          6360 => x"fe119013",
          6361 => x"08595658",
          6362 => x"55757426",
          6363 => x"9138757c",
          6364 => x"0c81e439",
          6365 => x"815b81cc",
          6366 => x"39825b81",
          6367 => x"c73981dc",
          6368 => x"cc087533",
          6369 => x"55597381",
          6370 => x"2e098106",
          6371 => x"bf388275",
          6372 => x"5f577652",
          6373 => x"923df005",
          6374 => x"51c1f43f",
          6375 => x"81dccc08",
          6376 => x"ff2ed138",
          6377 => x"81dccc08",
          6378 => x"812ece38",
          6379 => x"81dccc08",
          6380 => x"307081dc",
          6381 => x"cc080780",
          6382 => x"257a0581",
          6383 => x"197f5359",
          6384 => x"5a549814",
          6385 => x"087726ca",
          6386 => x"3880f939",
          6387 => x"a4150881",
          6388 => x"dccc0857",
          6389 => x"58759838",
          6390 => x"77528118",
          6391 => x"7d5258ff",
          6392 => x"bf8d3f81",
          6393 => x"dccc085b",
          6394 => x"81dccc08",
          6395 => x"80d6387c",
          6396 => x"70337712",
          6397 => x"ff1a5d52",
          6398 => x"56547482",
          6399 => x"2e098106",
          6400 => x"9e38b414",
          6401 => x"51ffbbcb",
          6402 => x"3f81dccc",
          6403 => x"0883ffff",
          6404 => x"06703070",
          6405 => x"80251b82",
          6406 => x"19595b51",
          6407 => x"549b39b4",
          6408 => x"1451ffbb",
          6409 => x"c53f81dc",
          6410 => x"cc08f00a",
          6411 => x"06703070",
          6412 => x"80251b84",
          6413 => x"19595b51",
          6414 => x"547583ff",
          6415 => x"067a5856",
          6416 => x"79ff9238",
          6417 => x"787c0c7c",
          6418 => x"7990120c",
          6419 => x"84113381",
          6420 => x"07565474",
          6421 => x"8415347a",
          6422 => x"81dccc0c",
          6423 => x"923d0d04",
          6424 => x"f93d0d79",
          6425 => x"8a3dfc05",
          6426 => x"53705257",
          6427 => x"e3dd3f81",
          6428 => x"dccc0856",
          6429 => x"81dccc08",
          6430 => x"81a83891",
          6431 => x"17335675",
          6432 => x"81a03890",
          6433 => x"17337081",
          6434 => x"2a708106",
          6435 => x"51555587",
          6436 => x"5573802e",
          6437 => x"818e3894",
          6438 => x"17085473",
          6439 => x"8c180827",
          6440 => x"81803873",
          6441 => x"9b3881dc",
          6442 => x"cc085388",
          6443 => x"17085276",
          6444 => x"51c48c3f",
          6445 => x"81dccc08",
          6446 => x"7488190c",
          6447 => x"5680c939",
          6448 => x"98170852",
          6449 => x"7651ffbf",
          6450 => x"c63f81dc",
          6451 => x"cc08ff2e",
          6452 => x"09810683",
          6453 => x"38815681",
          6454 => x"dccc0881",
          6455 => x"2e098106",
          6456 => x"85388256",
          6457 => x"a33975a0",
          6458 => x"38775481",
          6459 => x"dccc0898",
          6460 => x"15082794",
          6461 => x"38981708",
          6462 => x"5381dccc",
          6463 => x"08527651",
          6464 => x"c3bd3f81",
          6465 => x"dccc0856",
          6466 => x"9417088c",
          6467 => x"180c9017",
          6468 => x"3380c007",
          6469 => x"54739018",
          6470 => x"3475802e",
          6471 => x"85387591",
          6472 => x"18347555",
          6473 => x"7481dccc",
          6474 => x"0c893d0d",
          6475 => x"04e23d0d",
          6476 => x"8253a03d",
          6477 => x"ffa40552",
          6478 => x"a13d51da",
          6479 => x"e43f81dc",
          6480 => x"cc085581",
          6481 => x"dccc0881",
          6482 => x"f5387845",
          6483 => x"a13d0852",
          6484 => x"953d7052",
          6485 => x"58d1ae3f",
          6486 => x"81dccc08",
          6487 => x"5581dccc",
          6488 => x"0881db38",
          6489 => x"0280fb05",
          6490 => x"3370852a",
          6491 => x"70810651",
          6492 => x"55568655",
          6493 => x"7381c738",
          6494 => x"75982b54",
          6495 => x"80742481",
          6496 => x"bd380280",
          6497 => x"d6053370",
          6498 => x"81065854",
          6499 => x"87557681",
          6500 => x"ad386b52",
          6501 => x"7851ccc5",
          6502 => x"3f81dccc",
          6503 => x"0874842a",
          6504 => x"70810651",
          6505 => x"55567380",
          6506 => x"2e80d438",
          6507 => x"785481dc",
          6508 => x"cc089415",
          6509 => x"082e8186",
          6510 => x"38735a81",
          6511 => x"dccc085c",
          6512 => x"76528a3d",
          6513 => x"705254c7",
          6514 => x"b53f81dc",
          6515 => x"cc085581",
          6516 => x"dccc0880",
          6517 => x"e93881dc",
          6518 => x"cc085273",
          6519 => x"51cce53f",
          6520 => x"81dccc08",
          6521 => x"5581dccc",
          6522 => x"08863887",
          6523 => x"5580cf39",
          6524 => x"81dccc08",
          6525 => x"842e8838",
          6526 => x"81dccc08",
          6527 => x"80c03877",
          6528 => x"51cec23f",
          6529 => x"81dccc08",
          6530 => x"81dccc08",
          6531 => x"307081dc",
          6532 => x"cc080780",
          6533 => x"25515555",
          6534 => x"75802e94",
          6535 => x"3873802e",
          6536 => x"8f388053",
          6537 => x"75527751",
          6538 => x"c1953f81",
          6539 => x"dccc0855",
          6540 => x"748c3878",
          6541 => x"51ffbafe",
          6542 => x"3f81dccc",
          6543 => x"08557481",
          6544 => x"dccc0ca0",
          6545 => x"3d0d04e9",
          6546 => x"3d0d8253",
          6547 => x"993dc005",
          6548 => x"529a3d51",
          6549 => x"d8cb3f81",
          6550 => x"dccc0854",
          6551 => x"81dccc08",
          6552 => x"82b03878",
          6553 => x"5e69528e",
          6554 => x"3d705258",
          6555 => x"cf973f81",
          6556 => x"dccc0854",
          6557 => x"81dccc08",
          6558 => x"86388854",
          6559 => x"82943981",
          6560 => x"dccc0884",
          6561 => x"2e098106",
          6562 => x"82883802",
          6563 => x"80df0533",
          6564 => x"70852a81",
          6565 => x"06515586",
          6566 => x"547481f6",
          6567 => x"38785a74",
          6568 => x"528a3d70",
          6569 => x"5257c1c3",
          6570 => x"3f81dccc",
          6571 => x"08755556",
          6572 => x"81dccc08",
          6573 => x"83388754",
          6574 => x"81dccc08",
          6575 => x"812e0981",
          6576 => x"06833882",
          6577 => x"5481dccc",
          6578 => x"08ff2e09",
          6579 => x"81068638",
          6580 => x"815481b4",
          6581 => x"397381b0",
          6582 => x"3881dccc",
          6583 => x"08527851",
          6584 => x"c4a43f81",
          6585 => x"dccc0854",
          6586 => x"81dccc08",
          6587 => x"819a388b",
          6588 => x"53a052b4",
          6589 => x"1951ffb7",
          6590 => x"8c3f7854",
          6591 => x"ae0bb415",
          6592 => x"34785490",
          6593 => x"0bbf1534",
          6594 => x"8288b20a",
          6595 => x"5280ca19",
          6596 => x"51ffb69f",
          6597 => x"3f755378",
          6598 => x"b4115351",
          6599 => x"c9f83fa0",
          6600 => x"5378b411",
          6601 => x"5380d405",
          6602 => x"51ffb6b6",
          6603 => x"3f7854ae",
          6604 => x"0b80d515",
          6605 => x"347f5378",
          6606 => x"80d41153",
          6607 => x"51c9d73f",
          6608 => x"7854810b",
          6609 => x"83153477",
          6610 => x"51cba43f",
          6611 => x"81dccc08",
          6612 => x"5481dccc",
          6613 => x"08b23882",
          6614 => x"88b20a52",
          6615 => x"64960551",
          6616 => x"ffb5d03f",
          6617 => x"75536452",
          6618 => x"7851c9aa",
          6619 => x"3f645490",
          6620 => x"0b8b1534",
          6621 => x"7854810b",
          6622 => x"83153478",
          6623 => x"51ffb8b6",
          6624 => x"3f81dccc",
          6625 => x"08548b39",
          6626 => x"80537552",
          6627 => x"7651ffbe",
          6628 => x"ae3f7381",
          6629 => x"dccc0c99",
          6630 => x"3d0d04da",
          6631 => x"3d0da93d",
          6632 => x"840551d2",
          6633 => x"f13f8253",
          6634 => x"a83dff84",
          6635 => x"0552a93d",
          6636 => x"51d5ee3f",
          6637 => x"81dccc08",
          6638 => x"5581dccc",
          6639 => x"0882d338",
          6640 => x"784da93d",
          6641 => x"08529d3d",
          6642 => x"705258cc",
          6643 => x"b83f81dc",
          6644 => x"cc085581",
          6645 => x"dccc0882",
          6646 => x"b9380281",
          6647 => x"9b053381",
          6648 => x"a0065486",
          6649 => x"557382aa",
          6650 => x"38a053a4",
          6651 => x"3d0852a8",
          6652 => x"3dff8805",
          6653 => x"51ffb4ea",
          6654 => x"3fac5377",
          6655 => x"52923d70",
          6656 => x"5254ffb4",
          6657 => x"dd3faa3d",
          6658 => x"08527351",
          6659 => x"cbf73f81",
          6660 => x"dccc0855",
          6661 => x"81dccc08",
          6662 => x"9538636f",
          6663 => x"2e098106",
          6664 => x"883865a2",
          6665 => x"3d082e92",
          6666 => x"38885581",
          6667 => x"e53981dc",
          6668 => x"cc08842e",
          6669 => x"09810681",
          6670 => x"b8387351",
          6671 => x"c9b13f81",
          6672 => x"dccc0855",
          6673 => x"81dccc08",
          6674 => x"81c83868",
          6675 => x"569353a8",
          6676 => x"3dff9505",
          6677 => x"528d1651",
          6678 => x"ffb4873f",
          6679 => x"02af0533",
          6680 => x"8b17348b",
          6681 => x"16337084",
          6682 => x"2a708106",
          6683 => x"51555573",
          6684 => x"893874a0",
          6685 => x"0754738b",
          6686 => x"17347854",
          6687 => x"810b8315",
          6688 => x"348b1633",
          6689 => x"70842a70",
          6690 => x"81065155",
          6691 => x"5573802e",
          6692 => x"80e5386e",
          6693 => x"642e80df",
          6694 => x"38755278",
          6695 => x"51c6be3f",
          6696 => x"81dccc08",
          6697 => x"527851ff",
          6698 => x"b7bb3f82",
          6699 => x"5581dccc",
          6700 => x"08802e80",
          6701 => x"dd3881dc",
          6702 => x"cc085278",
          6703 => x"51ffb5af",
          6704 => x"3f81dccc",
          6705 => x"087980d4",
          6706 => x"11585855",
          6707 => x"81dccc08",
          6708 => x"80c03881",
          6709 => x"16335473",
          6710 => x"ae2e0981",
          6711 => x"06993863",
          6712 => x"53755276",
          6713 => x"51c6af3f",
          6714 => x"7854810b",
          6715 => x"83153487",
          6716 => x"3981dccc",
          6717 => x"089c3877",
          6718 => x"51c8ca3f",
          6719 => x"81dccc08",
          6720 => x"5581dccc",
          6721 => x"088c3878",
          6722 => x"51ffb5aa",
          6723 => x"3f81dccc",
          6724 => x"08557481",
          6725 => x"dccc0ca8",
          6726 => x"3d0d04ed",
          6727 => x"3d0d0280",
          6728 => x"db053302",
          6729 => x"840580df",
          6730 => x"05335757",
          6731 => x"8253953d",
          6732 => x"d0055296",
          6733 => x"3d51d2e9",
          6734 => x"3f81dccc",
          6735 => x"085581dc",
          6736 => x"cc0880cf",
          6737 => x"38785a65",
          6738 => x"52953dd4",
          6739 => x"0551c9b5",
          6740 => x"3f81dccc",
          6741 => x"085581dc",
          6742 => x"cc08b838",
          6743 => x"0280cf05",
          6744 => x"3381a006",
          6745 => x"54865573",
          6746 => x"aa3875a7",
          6747 => x"06617109",
          6748 => x"8b123371",
          6749 => x"067a7406",
          6750 => x"07515755",
          6751 => x"56748b15",
          6752 => x"34785481",
          6753 => x"0b831534",
          6754 => x"7851ffb4",
          6755 => x"a93f81dc",
          6756 => x"cc085574",
          6757 => x"81dccc0c",
          6758 => x"953d0d04",
          6759 => x"ef3d0d64",
          6760 => x"56825393",
          6761 => x"3dd00552",
          6762 => x"943d51d1",
          6763 => x"f43f81dc",
          6764 => x"cc085581",
          6765 => x"dccc0880",
          6766 => x"cb387658",
          6767 => x"6352933d",
          6768 => x"d40551c8",
          6769 => x"c03f81dc",
          6770 => x"cc085581",
          6771 => x"dccc08b4",
          6772 => x"380280c7",
          6773 => x"053381a0",
          6774 => x"06548655",
          6775 => x"73a63884",
          6776 => x"16228617",
          6777 => x"2271902b",
          6778 => x"07535496",
          6779 => x"1f51ffb0",
          6780 => x"c23f7654",
          6781 => x"810b8315",
          6782 => x"347651ff",
          6783 => x"b3b83f81",
          6784 => x"dccc0855",
          6785 => x"7481dccc",
          6786 => x"0c933d0d",
          6787 => x"04ea3d0d",
          6788 => x"696b5c5a",
          6789 => x"8053983d",
          6790 => x"d0055299",
          6791 => x"3d51d181",
          6792 => x"3f81dccc",
          6793 => x"0881dccc",
          6794 => x"08307081",
          6795 => x"dccc0807",
          6796 => x"80255155",
          6797 => x"5779802e",
          6798 => x"81853881",
          6799 => x"70750655",
          6800 => x"5573802e",
          6801 => x"80f9387b",
          6802 => x"5d805f80",
          6803 => x"528d3d70",
          6804 => x"5254ffbe",
          6805 => x"a93f81dc",
          6806 => x"cc085781",
          6807 => x"dccc0880",
          6808 => x"d1387452",
          6809 => x"7351c3dc",
          6810 => x"3f81dccc",
          6811 => x"085781dc",
          6812 => x"cc08bf38",
          6813 => x"81dccc08",
          6814 => x"81dccc08",
          6815 => x"655b5956",
          6816 => x"78188119",
          6817 => x"7b185659",
          6818 => x"55743374",
          6819 => x"34811656",
          6820 => x"8a7827ec",
          6821 => x"388b5675",
          6822 => x"1a548074",
          6823 => x"3475802e",
          6824 => x"9e38ff16",
          6825 => x"701b7033",
          6826 => x"51555673",
          6827 => x"a02ee838",
          6828 => x"8e397684",
          6829 => x"2e098106",
          6830 => x"8638807a",
          6831 => x"34805776",
          6832 => x"30707807",
          6833 => x"80255154",
          6834 => x"7a802e80",
          6835 => x"c1387380",
          6836 => x"2ebc387b",
          6837 => x"a0110853",
          6838 => x"51ffb193",
          6839 => x"3f81dccc",
          6840 => x"085781dc",
          6841 => x"cc08a738",
          6842 => x"7b703355",
          6843 => x"5580c356",
          6844 => x"73832e8b",
          6845 => x"3880e456",
          6846 => x"73842e83",
          6847 => x"38a75675",
          6848 => x"15b40551",
          6849 => x"ffade33f",
          6850 => x"81dccc08",
          6851 => x"7b0c7681",
          6852 => x"dccc0c98",
          6853 => x"3d0d04e6",
          6854 => x"3d0d8253",
          6855 => x"9c3dffb8",
          6856 => x"05529d3d",
          6857 => x"51cefa3f",
          6858 => x"81dccc08",
          6859 => x"81dccc08",
          6860 => x"565481dc",
          6861 => x"cc088398",
          6862 => x"388b53a0",
          6863 => x"528b3d70",
          6864 => x"5259ffae",
          6865 => x"c03f736d",
          6866 => x"70337081",
          6867 => x"ff065257",
          6868 => x"55579f74",
          6869 => x"2781bc38",
          6870 => x"78587481",
          6871 => x"ff066d81",
          6872 => x"054e7052",
          6873 => x"55ffaf89",
          6874 => x"3f81dccc",
          6875 => x"08802ea5",
          6876 => x"386c7033",
          6877 => x"70535754",
          6878 => x"ffaefd3f",
          6879 => x"81dccc08",
          6880 => x"802e8d38",
          6881 => x"74882b76",
          6882 => x"076d8105",
          6883 => x"4e558639",
          6884 => x"81dccc08",
          6885 => x"55ff9f15",
          6886 => x"7083ffff",
          6887 => x"06515473",
          6888 => x"99268a38",
          6889 => x"e0157083",
          6890 => x"ffff0656",
          6891 => x"5480ff75",
          6892 => x"27873881",
          6893 => x"cb9c1533",
          6894 => x"5574802e",
          6895 => x"a3387452",
          6896 => x"81cd9c51",
          6897 => x"ffae893f",
          6898 => x"81dccc08",
          6899 => x"933881ff",
          6900 => x"75278838",
          6901 => x"76892688",
          6902 => x"388b398a",
          6903 => x"77278638",
          6904 => x"865581ec",
          6905 => x"3981ff75",
          6906 => x"278f3874",
          6907 => x"882a5473",
          6908 => x"78708105",
          6909 => x"5a348117",
          6910 => x"57747870",
          6911 => x"81055a34",
          6912 => x"81176d70",
          6913 => x"337081ff",
          6914 => x"06525755",
          6915 => x"57739f26",
          6916 => x"fec8388b",
          6917 => x"3d335486",
          6918 => x"557381e5",
          6919 => x"2e81b138",
          6920 => x"76802e99",
          6921 => x"3802a705",
          6922 => x"55761570",
          6923 => x"33515473",
          6924 => x"a02e0981",
          6925 => x"068738ff",
          6926 => x"175776ed",
          6927 => x"38794180",
          6928 => x"43805291",
          6929 => x"3d705255",
          6930 => x"ffbab33f",
          6931 => x"81dccc08",
          6932 => x"5481dccc",
          6933 => x"0880f738",
          6934 => x"81527451",
          6935 => x"ffbfe53f",
          6936 => x"81dccc08",
          6937 => x"5481dccc",
          6938 => x"088d3876",
          6939 => x"80c43867",
          6940 => x"54e57434",
          6941 => x"80c63981",
          6942 => x"dccc0884",
          6943 => x"2e098106",
          6944 => x"80cc3880",
          6945 => x"5476742e",
          6946 => x"80c43881",
          6947 => x"527451ff",
          6948 => x"bdb03f81",
          6949 => x"dccc0854",
          6950 => x"81dccc08",
          6951 => x"b138a053",
          6952 => x"81dccc08",
          6953 => x"526751ff",
          6954 => x"abdb3f67",
          6955 => x"54880b8b",
          6956 => x"15348b53",
          6957 => x"78526751",
          6958 => x"ffaba73f",
          6959 => x"7954810b",
          6960 => x"83153479",
          6961 => x"51ffadee",
          6962 => x"3f81dccc",
          6963 => x"08547355",
          6964 => x"7481dccc",
          6965 => x"0c9c3d0d",
          6966 => x"04f23d0d",
          6967 => x"60620288",
          6968 => x"0580cb05",
          6969 => x"33933dfc",
          6970 => x"05557254",
          6971 => x"405e5ad2",
          6972 => x"da3f81dc",
          6973 => x"cc085881",
          6974 => x"dccc0882",
          6975 => x"bd38911a",
          6976 => x"33587782",
          6977 => x"b5387c80",
          6978 => x"2e97388c",
          6979 => x"1a085978",
          6980 => x"9038901a",
          6981 => x"3370812a",
          6982 => x"70810651",
          6983 => x"55557390",
          6984 => x"38875482",
          6985 => x"97398258",
          6986 => x"82903981",
          6987 => x"58828b39",
          6988 => x"7e8a1122",
          6989 => x"70892b70",
          6990 => x"557f5456",
          6991 => x"5656fefc",
          6992 => x"b83fff14",
          6993 => x"7d067030",
          6994 => x"7072079f",
          6995 => x"2a81dccc",
          6996 => x"08058c19",
          6997 => x"087c405a",
          6998 => x"5d555581",
          6999 => x"77278838",
          7000 => x"98160877",
          7001 => x"26833882",
          7002 => x"57767756",
          7003 => x"59805674",
          7004 => x"527951ff",
          7005 => x"ae993f81",
          7006 => x"157f5555",
          7007 => x"98140875",
          7008 => x"26833882",
          7009 => x"5581dccc",
          7010 => x"08812eff",
          7011 => x"993881dc",
          7012 => x"cc08ff2e",
          7013 => x"ff953881",
          7014 => x"dccc088e",
          7015 => x"38811656",
          7016 => x"757b2e09",
          7017 => x"81068738",
          7018 => x"93397459",
          7019 => x"80567477",
          7020 => x"2e098106",
          7021 => x"ffb93887",
          7022 => x"5880ff39",
          7023 => x"7d802eba",
          7024 => x"38787b55",
          7025 => x"557a802e",
          7026 => x"b4388115",
          7027 => x"5673812e",
          7028 => x"09810683",
          7029 => x"38ff5675",
          7030 => x"5374527e",
          7031 => x"51ffafa8",
          7032 => x"3f81dccc",
          7033 => x"085881dc",
          7034 => x"cc0880ce",
          7035 => x"38748116",
          7036 => x"ff165656",
          7037 => x"5c73d338",
          7038 => x"8439ff19",
          7039 => x"5c7e7c8c",
          7040 => x"120c557d",
          7041 => x"802eb338",
          7042 => x"78881b0c",
          7043 => x"7c8c1b0c",
          7044 => x"901a3380",
          7045 => x"c0075473",
          7046 => x"901b3498",
          7047 => x"1508fe05",
          7048 => x"90160857",
          7049 => x"54757426",
          7050 => x"9138757b",
          7051 => x"3190160c",
          7052 => x"84153381",
          7053 => x"07547384",
          7054 => x"16347754",
          7055 => x"7381dccc",
          7056 => x"0c903d0d",
          7057 => x"04e93d0d",
          7058 => x"6b6d0288",
          7059 => x"0580eb05",
          7060 => x"339d3d54",
          7061 => x"5a5c59c5",
          7062 => x"bd3f8b56",
          7063 => x"800b81dc",
          7064 => x"cc08248b",
          7065 => x"f83881dc",
          7066 => x"cc088429",
          7067 => x"81dce805",
          7068 => x"70085155",
          7069 => x"74802e84",
          7070 => x"38807534",
          7071 => x"81dccc08",
          7072 => x"81ff065f",
          7073 => x"81527e51",
          7074 => x"ffa0d03f",
          7075 => x"81dccc08",
          7076 => x"81ff0670",
          7077 => x"81065657",
          7078 => x"8356748b",
          7079 => x"c0387682",
          7080 => x"2a708106",
          7081 => x"51558a56",
          7082 => x"748bb238",
          7083 => x"993dfc05",
          7084 => x"5383527e",
          7085 => x"51ffa4f0",
          7086 => x"3f81dccc",
          7087 => x"08993867",
          7088 => x"5574802e",
          7089 => x"92387482",
          7090 => x"8080268b",
          7091 => x"38ff1575",
          7092 => x"06557480",
          7093 => x"2e833881",
          7094 => x"4878802e",
          7095 => x"87388480",
          7096 => x"79269238",
          7097 => x"7881800a",
          7098 => x"268b38ff",
          7099 => x"19790655",
          7100 => x"74802e86",
          7101 => x"3893568a",
          7102 => x"e4397889",
          7103 => x"2a6e892a",
          7104 => x"70892b77",
          7105 => x"59484359",
          7106 => x"7a833881",
          7107 => x"56613070",
          7108 => x"80257707",
          7109 => x"51559156",
          7110 => x"748ac238",
          7111 => x"993df805",
          7112 => x"5381527e",
          7113 => x"51ffa480",
          7114 => x"3f815681",
          7115 => x"dccc088a",
          7116 => x"ac387783",
          7117 => x"2a707706",
          7118 => x"81dccc08",
          7119 => x"43564574",
          7120 => x"8338bf41",
          7121 => x"66558e56",
          7122 => x"6075268a",
          7123 => x"90387461",
          7124 => x"31704855",
          7125 => x"80ff7527",
          7126 => x"8a833893",
          7127 => x"56788180",
          7128 => x"2689fa38",
          7129 => x"77812a70",
          7130 => x"81065643",
          7131 => x"74802e95",
          7132 => x"38778706",
          7133 => x"5574822e",
          7134 => x"838d3877",
          7135 => x"81065574",
          7136 => x"802e8383",
          7137 => x"38778106",
          7138 => x"55935682",
          7139 => x"5e74802e",
          7140 => x"89cb3878",
          7141 => x"5a7d832e",
          7142 => x"09810680",
          7143 => x"e13878ae",
          7144 => x"3866912a",
          7145 => x"57810b81",
          7146 => x"cdc02256",
          7147 => x"5a74802e",
          7148 => x"9d387477",
          7149 => x"26983881",
          7150 => x"cdc05679",
          7151 => x"10821770",
          7152 => x"2257575a",
          7153 => x"74802e86",
          7154 => x"38767527",
          7155 => x"ee387952",
          7156 => x"6651fef7",
          7157 => x"a43f81dc",
          7158 => x"cc088429",
          7159 => x"84870570",
          7160 => x"892a5e55",
          7161 => x"a05c800b",
          7162 => x"81dccc08",
          7163 => x"fc808a05",
          7164 => x"5644fdff",
          7165 => x"f00a7527",
          7166 => x"80ec3888",
          7167 => x"d33978ae",
          7168 => x"38668c2a",
          7169 => x"57810b81",
          7170 => x"cdb02256",
          7171 => x"5a74802e",
          7172 => x"9d387477",
          7173 => x"26983881",
          7174 => x"cdb05679",
          7175 => x"10821770",
          7176 => x"2257575a",
          7177 => x"74802e86",
          7178 => x"38767527",
          7179 => x"ee387952",
          7180 => x"6651fef6",
          7181 => x"c43f81dc",
          7182 => x"cc081084",
          7183 => x"055781dc",
          7184 => x"cc089ff5",
          7185 => x"26963881",
          7186 => x"0b81dccc",
          7187 => x"081081dc",
          7188 => x"cc080571",
          7189 => x"11722a83",
          7190 => x"0559565e",
          7191 => x"83ff1789",
          7192 => x"2a5d815c",
          7193 => x"a044601c",
          7194 => x"7d116505",
          7195 => x"697012ff",
          7196 => x"05713070",
          7197 => x"72067431",
          7198 => x"5c525957",
          7199 => x"59407d83",
          7200 => x"2e098106",
          7201 => x"8938761c",
          7202 => x"6018415c",
          7203 => x"8439761d",
          7204 => x"5d799029",
          7205 => x"18706231",
          7206 => x"68585155",
          7207 => x"74762687",
          7208 => x"af38757c",
          7209 => x"317d317a",
          7210 => x"53706531",
          7211 => x"5255fef5",
          7212 => x"c83f81dc",
          7213 => x"cc08587d",
          7214 => x"832e0981",
          7215 => x"069b3881",
          7216 => x"dccc0883",
          7217 => x"fff52680",
          7218 => x"dd387887",
          7219 => x"83387981",
          7220 => x"2a5978fd",
          7221 => x"be3886f8",
          7222 => x"397d822e",
          7223 => x"09810680",
          7224 => x"c53883ff",
          7225 => x"f50b81dc",
          7226 => x"cc0827a0",
          7227 => x"38788f38",
          7228 => x"791a5574",
          7229 => x"80c02686",
          7230 => x"387459fd",
          7231 => x"96396281",
          7232 => x"06557480",
          7233 => x"2e8f3883",
          7234 => x"5efd8839",
          7235 => x"81dccc08",
          7236 => x"9ff52692",
          7237 => x"387886b8",
          7238 => x"38791a59",
          7239 => x"81807927",
          7240 => x"fcf13886",
          7241 => x"ab398055",
          7242 => x"7d812e09",
          7243 => x"81068338",
          7244 => x"7d559ff5",
          7245 => x"78278b38",
          7246 => x"74810655",
          7247 => x"8e567486",
          7248 => x"9c388480",
          7249 => x"5380527a",
          7250 => x"51ffa2b9",
          7251 => x"3f8b5381",
          7252 => x"cbd8527a",
          7253 => x"51ffa28a",
          7254 => x"3f848052",
          7255 => x"8b1b51ff",
          7256 => x"a1b33f79",
          7257 => x"8d1c347b",
          7258 => x"83ffff06",
          7259 => x"528e1b51",
          7260 => x"ffa1a23f",
          7261 => x"810b901c",
          7262 => x"347d8332",
          7263 => x"70307096",
          7264 => x"2a848006",
          7265 => x"54515591",
          7266 => x"1b51ffa1",
          7267 => x"883f6655",
          7268 => x"7483ffff",
          7269 => x"26903874",
          7270 => x"83ffff06",
          7271 => x"52931b51",
          7272 => x"ffa0f23f",
          7273 => x"8a397452",
          7274 => x"a01b51ff",
          7275 => x"a1853ff8",
          7276 => x"0b951c34",
          7277 => x"bf52981b",
          7278 => x"51ffa0d9",
          7279 => x"3f81ff52",
          7280 => x"9a1b51ff",
          7281 => x"a0cf3f60",
          7282 => x"529c1b51",
          7283 => x"ffa0e43f",
          7284 => x"7d832e09",
          7285 => x"810680cb",
          7286 => x"388288b2",
          7287 => x"0a5280c3",
          7288 => x"1b51ffa0",
          7289 => x"ce3f7c52",
          7290 => x"a41b51ff",
          7291 => x"a0c53f82",
          7292 => x"52ac1b51",
          7293 => x"ffa0bc3f",
          7294 => x"8152b01b",
          7295 => x"51ffa095",
          7296 => x"3f8652b2",
          7297 => x"1b51ffa0",
          7298 => x"8c3fff80",
          7299 => x"0b80c01c",
          7300 => x"34a90b80",
          7301 => x"c21c3493",
          7302 => x"5381cbe4",
          7303 => x"5280c71b",
          7304 => x"51ae3982",
          7305 => x"88b20a52",
          7306 => x"a71b51ff",
          7307 => x"a0853f7c",
          7308 => x"83ffff06",
          7309 => x"52961b51",
          7310 => x"ff9fda3f",
          7311 => x"ff800ba4",
          7312 => x"1c34a90b",
          7313 => x"a61c3493",
          7314 => x"5381cbf8",
          7315 => x"52ab1b51",
          7316 => x"ffa08f3f",
          7317 => x"82d4d552",
          7318 => x"83fe1b70",
          7319 => x"5259ff9f",
          7320 => x"b43f8154",
          7321 => x"60537a52",
          7322 => x"7e51ff9b",
          7323 => x"d73f8156",
          7324 => x"81dccc08",
          7325 => x"83e7387d",
          7326 => x"832e0981",
          7327 => x"0680ee38",
          7328 => x"75546086",
          7329 => x"05537a52",
          7330 => x"7e51ff9b",
          7331 => x"b73f8480",
          7332 => x"5380527a",
          7333 => x"51ff9fed",
          7334 => x"3f848b85",
          7335 => x"a4d2527a",
          7336 => x"51ff9f8f",
          7337 => x"3f868a85",
          7338 => x"e4f25283",
          7339 => x"e41b51ff",
          7340 => x"9f813fff",
          7341 => x"185283e8",
          7342 => x"1b51ff9e",
          7343 => x"f63f8252",
          7344 => x"83ec1b51",
          7345 => x"ff9eec3f",
          7346 => x"82d4d552",
          7347 => x"7851ff9e",
          7348 => x"c43f7554",
          7349 => x"60870553",
          7350 => x"7a527e51",
          7351 => x"ff9ae53f",
          7352 => x"75546016",
          7353 => x"537a527e",
          7354 => x"51ff9ad8",
          7355 => x"3f655380",
          7356 => x"527a51ff",
          7357 => x"9f8f3f7f",
          7358 => x"5680587d",
          7359 => x"832e0981",
          7360 => x"069a38f8",
          7361 => x"527a51ff",
          7362 => x"9ea93fff",
          7363 => x"52841b51",
          7364 => x"ff9ea03f",
          7365 => x"f00a5288",
          7366 => x"1b519139",
          7367 => x"87fffff8",
          7368 => x"557d812e",
          7369 => x"8338f855",
          7370 => x"74527a51",
          7371 => x"ff9e843f",
          7372 => x"7c556157",
          7373 => x"74622683",
          7374 => x"38745776",
          7375 => x"5475537a",
          7376 => x"527e51ff",
          7377 => x"99fe3f81",
          7378 => x"dccc0882",
          7379 => x"87388480",
          7380 => x"5381dccc",
          7381 => x"08527a51",
          7382 => x"ff9eaa3f",
          7383 => x"76167578",
          7384 => x"31565674",
          7385 => x"cd388118",
          7386 => x"5877802e",
          7387 => x"ff8d3879",
          7388 => x"557d832e",
          7389 => x"83386355",
          7390 => x"61577462",
          7391 => x"26833874",
          7392 => x"57765475",
          7393 => x"537a527e",
          7394 => x"51ff99b8",
          7395 => x"3f81dccc",
          7396 => x"0881c138",
          7397 => x"76167578",
          7398 => x"31565674",
          7399 => x"db388c56",
          7400 => x"7d832e93",
          7401 => x"38865666",
          7402 => x"83ffff26",
          7403 => x"8a388456",
          7404 => x"7d822e83",
          7405 => x"38815664",
          7406 => x"81065877",
          7407 => x"80fe3884",
          7408 => x"80537752",
          7409 => x"7a51ff9d",
          7410 => x"bc3f82d4",
          7411 => x"d5527851",
          7412 => x"ff9cc23f",
          7413 => x"83be1b55",
          7414 => x"77753481",
          7415 => x"0b811634",
          7416 => x"810b8216",
          7417 => x"34778316",
          7418 => x"34758416",
          7419 => x"34606705",
          7420 => x"5680fdc1",
          7421 => x"527551fe",
          7422 => x"eeff3ffe",
          7423 => x"0b851634",
          7424 => x"81dccc08",
          7425 => x"822abf07",
          7426 => x"56758616",
          7427 => x"3481dccc",
          7428 => x"08871634",
          7429 => x"605283c6",
          7430 => x"1b51ff9c",
          7431 => x"963f6652",
          7432 => x"83ca1b51",
          7433 => x"ff9c8c3f",
          7434 => x"81547753",
          7435 => x"7a527e51",
          7436 => x"ff98913f",
          7437 => x"815681dc",
          7438 => x"cc08a238",
          7439 => x"80538052",
          7440 => x"7e51ff99",
          7441 => x"e33f8156",
          7442 => x"81dccc08",
          7443 => x"90388939",
          7444 => x"8e568a39",
          7445 => x"81568639",
          7446 => x"81dccc08",
          7447 => x"567581dc",
          7448 => x"cc0c993d",
          7449 => x"0d04f53d",
          7450 => x"0d7d605b",
          7451 => x"59807960",
          7452 => x"ff055a57",
          7453 => x"57767825",
          7454 => x"b4388d3d",
          7455 => x"f8115555",
          7456 => x"8153fc15",
          7457 => x"527951c9",
          7458 => x"dc3f7a81",
          7459 => x"2e098106",
          7460 => x"9c388c3d",
          7461 => x"3355748d",
          7462 => x"2edb3874",
          7463 => x"76708105",
          7464 => x"58348117",
          7465 => x"57748a2e",
          7466 => x"098106c9",
          7467 => x"38807634",
          7468 => x"78557683",
          7469 => x"38765574",
          7470 => x"81dccc0c",
          7471 => x"8d3d0d04",
          7472 => x"fa3d0d78",
          7473 => x"70087055",
          7474 => x"56577480",
          7475 => x"2e80ea38",
          7476 => x"8e397477",
          7477 => x"0c851433",
          7478 => x"5380de39",
          7479 => x"81155580",
          7480 => x"75335556",
          7481 => x"73a02e83",
          7482 => x"38815673",
          7483 => x"30709f2a",
          7484 => x"77065153",
          7485 => x"72e63873",
          7486 => x"a02e0981",
          7487 => x"06883872",
          7488 => x"75708105",
          7489 => x"57347256",
          7490 => x"75902981",
          7491 => x"d9dc0577",
          7492 => x"08537008",
          7493 => x"5254fef3",
          7494 => x"f83f81dc",
          7495 => x"cc088b38",
          7496 => x"84143353",
          7497 => x"72812eff",
          7498 => x"a9388116",
          7499 => x"7081ff06",
          7500 => x"57539676",
          7501 => x"27d238ff",
          7502 => x"537281dc",
          7503 => x"cc0c883d",
          7504 => x"0d04ff3d",
          7505 => x"0d735271",
          7506 => x"9326818e",
          7507 => x"38718429",
          7508 => x"81c4fc05",
          7509 => x"52710804",
          7510 => x"81cee851",
          7511 => x"81803981",
          7512 => x"cef45180",
          7513 => x"f93981cf",
          7514 => x"885180f2",
          7515 => x"3981cf9c",
          7516 => x"5180eb39",
          7517 => x"81cfac51",
          7518 => x"80e43981",
          7519 => x"cfbc5180",
          7520 => x"dd3981cf",
          7521 => x"d05180d6",
          7522 => x"3981cfe0",
          7523 => x"5180cf39",
          7524 => x"81cff851",
          7525 => x"80c83981",
          7526 => x"d0905180",
          7527 => x"c13981d0",
          7528 => x"a851bb39",
          7529 => x"81d0c451",
          7530 => x"b53981d0",
          7531 => x"d851af39",
          7532 => x"81d18451",
          7533 => x"a93981d1",
          7534 => x"9851a339",
          7535 => x"81d1b851",
          7536 => x"9d3981d1",
          7537 => x"cc519739",
          7538 => x"81d1e451",
          7539 => x"913981d1",
          7540 => x"fc518b39",
          7541 => x"81d29451",
          7542 => x"853981d2",
          7543 => x"a051ff86",
          7544 => x"9f3f833d",
          7545 => x"0d04fb3d",
          7546 => x"0d777956",
          7547 => x"567487e7",
          7548 => x"268a3874",
          7549 => x"527587e8",
          7550 => x"29519139",
          7551 => x"87e85274",
          7552 => x"51feeaf5",
          7553 => x"3f81dccc",
          7554 => x"08527551",
          7555 => x"feeaea3f",
          7556 => x"81dccc08",
          7557 => x"54795375",
          7558 => x"5281d2b0",
          7559 => x"51ff8bc4",
          7560 => x"3f873d0d",
          7561 => x"04ec3d0d",
          7562 => x"66028405",
          7563 => x"80e30533",
          7564 => x"5b578068",
          7565 => x"7830707a",
          7566 => x"07732551",
          7567 => x"57595978",
          7568 => x"567787ff",
          7569 => x"26833881",
          7570 => x"56747607",
          7571 => x"7081ff06",
          7572 => x"51559356",
          7573 => x"7480ff38",
          7574 => x"81537652",
          7575 => x"8c3d7052",
          7576 => x"56c19d3f",
          7577 => x"81dccc08",
          7578 => x"5781dccc",
          7579 => x"08b83881",
          7580 => x"dccc0887",
          7581 => x"c098880c",
          7582 => x"81dccc08",
          7583 => x"59963dd4",
          7584 => x"05548480",
          7585 => x"53775275",
          7586 => x"51c5da3f",
          7587 => x"81dccc08",
          7588 => x"5781dccc",
          7589 => x"0890387a",
          7590 => x"5574802e",
          7591 => x"89387419",
          7592 => x"75195959",
          7593 => x"d839963d",
          7594 => x"d80551cd",
          7595 => x"c43f7630",
          7596 => x"70780780",
          7597 => x"257b3070",
          7598 => x"9f2a7206",
          7599 => x"51575156",
          7600 => x"74802e90",
          7601 => x"3881d2d4",
          7602 => x"5387c098",
          7603 => x"88085278",
          7604 => x"51fe933f",
          7605 => x"76567581",
          7606 => x"dccc0c96",
          7607 => x"3d0d04f9",
          7608 => x"3d0d7b02",
          7609 => x"8405b305",
          7610 => x"335758ff",
          7611 => x"5780537a",
          7612 => x"527951fe",
          7613 => x"b03f81dc",
          7614 => x"cc08a438",
          7615 => x"75802e88",
          7616 => x"3875812e",
          7617 => x"98389839",
          7618 => x"60557f54",
          7619 => x"81dccc53",
          7620 => x"7e527d51",
          7621 => x"772d81dc",
          7622 => x"cc085783",
          7623 => x"39770476",
          7624 => x"81dccc0c",
          7625 => x"893d0d04",
          7626 => x"f33d0d7f",
          7627 => x"6163028c",
          7628 => x"0580cf05",
          7629 => x"33737315",
          7630 => x"68415f5c",
          7631 => x"5c5e5e5e",
          7632 => x"7a5281d2",
          7633 => x"dc51ff89",
          7634 => x"9b3f81d2",
          7635 => x"e451ff83",
          7636 => x"af3f8055",
          7637 => x"74792780",
          7638 => x"fc387b90",
          7639 => x"2e89387b",
          7640 => x"a02ea738",
          7641 => x"80c63974",
          7642 => x"1853727a",
          7643 => x"278e3872",
          7644 => x"225281d2",
          7645 => x"e851ff88",
          7646 => x"eb3f8939",
          7647 => x"81d2f451",
          7648 => x"ff82fd3f",
          7649 => x"82155580",
          7650 => x"c3397418",
          7651 => x"53727a27",
          7652 => x"8e387208",
          7653 => x"5281d2dc",
          7654 => x"51ff88c8",
          7655 => x"3f893981",
          7656 => x"d2f051ff",
          7657 => x"82da3f84",
          7658 => x"1555a139",
          7659 => x"74185372",
          7660 => x"7a278e38",
          7661 => x"72335281",
          7662 => x"d2fc51ff",
          7663 => x"88a63f89",
          7664 => x"3981d384",
          7665 => x"51ff82b8",
          7666 => x"3f811555",
          7667 => x"a051ff81",
          7668 => x"d23fff80",
          7669 => x"3981d388",
          7670 => x"51ff82a4",
          7671 => x"3f805574",
          7672 => x"7927bc38",
          7673 => x"74187033",
          7674 => x"55538056",
          7675 => x"727a2783",
          7676 => x"38815680",
          7677 => x"539f7427",
          7678 => x"83388153",
          7679 => x"75730670",
          7680 => x"81ff0651",
          7681 => x"5372802e",
          7682 => x"8b387380",
          7683 => x"fe268538",
          7684 => x"73518339",
          7685 => x"a051ff81",
          7686 => x"8a3f8115",
          7687 => x"55c13981",
          7688 => x"d38c51ff",
          7689 => x"81da3f78",
          7690 => x"18791c5c",
          7691 => x"58fef6de",
          7692 => x"3f81dccc",
          7693 => x"08982b70",
          7694 => x"982c5157",
          7695 => x"76a02e09",
          7696 => x"8106ab38",
          7697 => x"fef6c73f",
          7698 => x"81dccc08",
          7699 => x"982b7098",
          7700 => x"2c70a032",
          7701 => x"7030729b",
          7702 => x"32703070",
          7703 => x"72077375",
          7704 => x"07065158",
          7705 => x"58595751",
          7706 => x"57807324",
          7707 => x"d738769b",
          7708 => x"2e098106",
          7709 => x"85388053",
          7710 => x"8c397c1e",
          7711 => x"53727826",
          7712 => x"fdbe38ff",
          7713 => x"537281dc",
          7714 => x"cc0c8f3d",
          7715 => x"0d04fc3d",
          7716 => x"0d029b05",
          7717 => x"3381d390",
          7718 => x"5381d394",
          7719 => x"5255ff86",
          7720 => x"c33f81d9",
          7721 => x"ac2251fe",
          7722 => x"ff9f3f81",
          7723 => x"d3a05481",
          7724 => x"d3ac5381",
          7725 => x"d9ad3352",
          7726 => x"81d3b451",
          7727 => x"ff86a53f",
          7728 => x"74802e85",
          7729 => x"38fefaea",
          7730 => x"3f863d0d",
          7731 => x"04fe3d0d",
          7732 => x"87c09680",
          7733 => x"0853feff",
          7734 => x"b83f8151",
          7735 => x"fef1c33f",
          7736 => x"81d3d051",
          7737 => x"fef3bb3f",
          7738 => x"8051fef1",
          7739 => x"b53f7281",
          7740 => x"2a708106",
          7741 => x"51527180",
          7742 => x"2e953881",
          7743 => x"51fef1a2",
          7744 => x"3f81d3e8",
          7745 => x"51fef39a",
          7746 => x"3f8051fe",
          7747 => x"f1943f72",
          7748 => x"822a7081",
          7749 => x"06515271",
          7750 => x"802e9538",
          7751 => x"8151fef1",
          7752 => x"813f81d3",
          7753 => x"fc51fef2",
          7754 => x"f93f8051",
          7755 => x"fef0f33f",
          7756 => x"72832a70",
          7757 => x"81065152",
          7758 => x"71802e95",
          7759 => x"388151fe",
          7760 => x"f0e03f81",
          7761 => x"d48c51fe",
          7762 => x"f2d83f80",
          7763 => x"51fef0d2",
          7764 => x"3f72842a",
          7765 => x"70810651",
          7766 => x"5271802e",
          7767 => x"95388151",
          7768 => x"fef0bf3f",
          7769 => x"81d4a051",
          7770 => x"fef2b73f",
          7771 => x"8051fef0",
          7772 => x"b13f7285",
          7773 => x"2a708106",
          7774 => x"51527180",
          7775 => x"2e953881",
          7776 => x"51fef09e",
          7777 => x"3f81d4b4",
          7778 => x"51fef296",
          7779 => x"3f8051fe",
          7780 => x"f0903f72",
          7781 => x"862a7081",
          7782 => x"06515271",
          7783 => x"802e9538",
          7784 => x"8151feef",
          7785 => x"fd3f81d4",
          7786 => x"c851fef1",
          7787 => x"f53f8051",
          7788 => x"feefef3f",
          7789 => x"72872a70",
          7790 => x"81065152",
          7791 => x"71802e95",
          7792 => x"388151fe",
          7793 => x"efdc3f81",
          7794 => x"d4dc51fe",
          7795 => x"f1d43f80",
          7796 => x"51feefce",
          7797 => x"3f72882a",
          7798 => x"70810651",
          7799 => x"5271802e",
          7800 => x"95388151",
          7801 => x"feefbb3f",
          7802 => x"81d4f051",
          7803 => x"fef1b33f",
          7804 => x"8051feef",
          7805 => x"ad3ffefd",
          7806 => x"a03f843d",
          7807 => x"0d04fb3d",
          7808 => x"0d777970",
          7809 => x"55565680",
          7810 => x"527551fe",
          7811 => x"e8f23f81",
          7812 => x"d9d83354",
          7813 => x"73a73881",
          7814 => x"5381d5b0",
          7815 => x"5281f3d0",
          7816 => x"51ffb9dc",
          7817 => x"3f81dccc",
          7818 => x"08307081",
          7819 => x"dccc0807",
          7820 => x"80258271",
          7821 => x"31515154",
          7822 => x"7381d9d8",
          7823 => x"3481d9d8",
          7824 => x"33547381",
          7825 => x"2e098106",
          7826 => x"ac3881f3",
          7827 => x"d0537452",
          7828 => x"7551f492",
          7829 => x"3f81dccc",
          7830 => x"08802e8c",
          7831 => x"3881dccc",
          7832 => x"0851fefd",
          7833 => x"9b3f8e39",
          7834 => x"81f3d051",
          7835 => x"c6833f82",
          7836 => x"0b81d9d8",
          7837 => x"3481d9d8",
          7838 => x"33547382",
          7839 => x"2e098106",
          7840 => x"89387452",
          7841 => x"7551ff83",
          7842 => x"b53f800b",
          7843 => x"81dccc0c",
          7844 => x"873d0d04",
          7845 => x"ce3d0d80",
          7846 => x"707181f3",
          7847 => x"cc0c5f5d",
          7848 => x"81527c51",
          7849 => x"ff88b43f",
          7850 => x"81dccc08",
          7851 => x"81ff0659",
          7852 => x"787d2e09",
          7853 => x"8106a238",
          7854 => x"81d5c052",
          7855 => x"963d7052",
          7856 => x"59ff82b6",
          7857 => x"3f7c5378",
          7858 => x"5281ddfc",
          7859 => x"51ffb7cf",
          7860 => x"3f81dccc",
          7861 => x"087d2e88",
          7862 => x"3881d5c4",
          7863 => x"518dc139",
          7864 => x"81705f5d",
          7865 => x"81d5fc51",
          7866 => x"fefc953f",
          7867 => x"963d7046",
          7868 => x"5a80f852",
          7869 => x"7951fe86",
          7870 => x"3fb43dff",
          7871 => x"840551f3",
          7872 => x"bf3f81dc",
          7873 => x"cc08902b",
          7874 => x"70902c51",
          7875 => x"597880c2",
          7876 => x"2e87b338",
          7877 => x"7880c224",
          7878 => x"b23878bd",
          7879 => x"2e81d538",
          7880 => x"78bd2490",
          7881 => x"3878802e",
          7882 => x"ffba3878",
          7883 => x"bc2e80da",
          7884 => x"388ae939",
          7885 => x"7880c02e",
          7886 => x"83a13878",
          7887 => x"80c02485",
          7888 => x"dd3878bf",
          7889 => x"2e829238",
          7890 => x"8ad23978",
          7891 => x"80f92e89",
          7892 => x"ea387880",
          7893 => x"f9249238",
          7894 => x"7880c32e",
          7895 => x"88983878",
          7896 => x"80f82e89",
          7897 => x"b1388ab4",
          7898 => x"39788183",
          7899 => x"2e8a9938",
          7900 => x"78818324",
          7901 => x"8b387881",
          7902 => x"822e89fd",
          7903 => x"388a9d39",
          7904 => x"7881852e",
          7905 => x"8a8f388a",
          7906 => x"9339b43d",
          7907 => x"ff801153",
          7908 => x"ff840551",
          7909 => x"ff82c23f",
          7910 => x"81dccc08",
          7911 => x"802efec4",
          7912 => x"38b43dfe",
          7913 => x"fc1153ff",
          7914 => x"840551ff",
          7915 => x"82ab3f81",
          7916 => x"dccc0880",
          7917 => x"2efead38",
          7918 => x"b43dfef8",
          7919 => x"1153ff84",
          7920 => x"0551ff82",
          7921 => x"943f81dc",
          7922 => x"cc088638",
          7923 => x"81dccc08",
          7924 => x"4281d680",
          7925 => x"51fefaa8",
          7926 => x"3f63635c",
          7927 => x"5a797b27",
          7928 => x"81f23861",
          7929 => x"59787a70",
          7930 => x"84055c0c",
          7931 => x"7a7a26f5",
          7932 => x"3881e139",
          7933 => x"b43dff80",
          7934 => x"1153ff84",
          7935 => x"0551ff81",
          7936 => x"d83f81dc",
          7937 => x"cc08802e",
          7938 => x"fdda38b4",
          7939 => x"3dfefc11",
          7940 => x"53ff8405",
          7941 => x"51ff81c1",
          7942 => x"3f81dccc",
          7943 => x"08802efd",
          7944 => x"c338b43d",
          7945 => x"fef81153",
          7946 => x"ff840551",
          7947 => x"ff81aa3f",
          7948 => x"81dccc08",
          7949 => x"802efdac",
          7950 => x"3881d690",
          7951 => x"51fef9c0",
          7952 => x"3f635a79",
          7953 => x"6327818c",
          7954 => x"38615979",
          7955 => x"7081055b",
          7956 => x"33793461",
          7957 => x"810542eb",
          7958 => x"39b43dff",
          7959 => x"801153ff",
          7960 => x"840551ff",
          7961 => x"80f33f81",
          7962 => x"dccc0880",
          7963 => x"2efcf538",
          7964 => x"b43dfefc",
          7965 => x"1153ff84",
          7966 => x"0551ff80",
          7967 => x"dc3f81dc",
          7968 => x"cc08802e",
          7969 => x"fcde38b4",
          7970 => x"3dfef811",
          7971 => x"53ff8405",
          7972 => x"51ff80c5",
          7973 => x"3f81dccc",
          7974 => x"08802efc",
          7975 => x"c73881d6",
          7976 => x"9c51fef8",
          7977 => x"db3f635a",
          7978 => x"796327a8",
          7979 => x"38617033",
          7980 => x"7b335e5a",
          7981 => x"5b787c2e",
          7982 => x"92387855",
          7983 => x"7a547933",
          7984 => x"53795281",
          7985 => x"d6ac51fe",
          7986 => x"fe9a3f81",
          7987 => x"1a628105",
          7988 => x"435ad539",
          7989 => x"81d6c451",
          7990 => x"82bd39b4",
          7991 => x"3dff8011",
          7992 => x"53ff8405",
          7993 => x"51fefff1",
          7994 => x"3f81dccc",
          7995 => x"0880df38",
          7996 => x"81d9c033",
          7997 => x"5978802e",
          7998 => x"893881d8",
          7999 => x"f8084480",
          8000 => x"cd3981d9",
          8001 => x"c1335978",
          8002 => x"802e8838",
          8003 => x"81d98008",
          8004 => x"44bc3981",
          8005 => x"d9c23359",
          8006 => x"78802e88",
          8007 => x"3881d988",
          8008 => x"0844ab39",
          8009 => x"81d9c333",
          8010 => x"5978802e",
          8011 => x"883881d9",
          8012 => x"9008449a",
          8013 => x"3981d9be",
          8014 => x"33597880",
          8015 => x"2e883881",
          8016 => x"d9980844",
          8017 => x"893981d9",
          8018 => x"a808fc80",
          8019 => x"0544b43d",
          8020 => x"fefc1153",
          8021 => x"ff840551",
          8022 => x"fefefe3f",
          8023 => x"81dccc08",
          8024 => x"80de3881",
          8025 => x"d9c03359",
          8026 => x"78802e89",
          8027 => x"3881d8fc",
          8028 => x"084380cc",
          8029 => x"3981d9c1",
          8030 => x"33597880",
          8031 => x"2e883881",
          8032 => x"d9840843",
          8033 => x"bb3981d9",
          8034 => x"c2335978",
          8035 => x"802e8838",
          8036 => x"81d98c08",
          8037 => x"43aa3981",
          8038 => x"d9c33359",
          8039 => x"78802e88",
          8040 => x"3881d994",
          8041 => x"08439939",
          8042 => x"81d9be33",
          8043 => x"5978802e",
          8044 => x"883881d9",
          8045 => x"9c084388",
          8046 => x"3981d9a8",
          8047 => x"08880543",
          8048 => x"b43dfef8",
          8049 => x"1153ff84",
          8050 => x"0551fefe",
          8051 => x"8c3f81dc",
          8052 => x"cc08802e",
          8053 => x"a7388062",
          8054 => x"5c5c7a88",
          8055 => x"2e833881",
          8056 => x"5c7a9032",
          8057 => x"70307072",
          8058 => x"079f2a70",
          8059 => x"7f065151",
          8060 => x"5a5a7880",
          8061 => x"2e88387a",
          8062 => x"a02e8338",
          8063 => x"884281d6",
          8064 => x"c851fef5",
          8065 => x"fb3fa055",
          8066 => x"63546153",
          8067 => x"62526351",
          8068 => x"f2963f81",
          8069 => x"d6d851fe",
          8070 => x"f5e63ff9",
          8071 => x"c739b43d",
          8072 => x"ff801153",
          8073 => x"ff840551",
          8074 => x"fefdae3f",
          8075 => x"81dccc08",
          8076 => x"802ef9b0",
          8077 => x"38b43dfe",
          8078 => x"fc1153ff",
          8079 => x"840551fe",
          8080 => x"fd973f81",
          8081 => x"dccc0880",
          8082 => x"2ea53863",
          8083 => x"590280cb",
          8084 => x"05337934",
          8085 => x"63810544",
          8086 => x"b43dfefc",
          8087 => x"1153ff84",
          8088 => x"0551fefc",
          8089 => x"f43f81dc",
          8090 => x"cc08e038",
          8091 => x"f8f63963",
          8092 => x"70335452",
          8093 => x"81d6e451",
          8094 => x"fefae93f",
          8095 => x"80f85279",
          8096 => x"51fefbba",
          8097 => x"3f794579",
          8098 => x"335978ae",
          8099 => x"2ef8d538",
          8100 => x"9f7927a0",
          8101 => x"38b43dfe",
          8102 => x"fc1153ff",
          8103 => x"840551fe",
          8104 => x"fcb73f81",
          8105 => x"dccc0880",
          8106 => x"2e913863",
          8107 => x"590280cb",
          8108 => x"05337934",
          8109 => x"63810544",
          8110 => x"ffb53981",
          8111 => x"d6f051fe",
          8112 => x"f4be3fff",
          8113 => x"aa39b43d",
          8114 => x"fef41153",
          8115 => x"ff840551",
          8116 => x"fefdf83f",
          8117 => x"81dccc08",
          8118 => x"802ef888",
          8119 => x"38b43dfe",
          8120 => x"f01153ff",
          8121 => x"840551fe",
          8122 => x"fde13f81",
          8123 => x"dccc0880",
          8124 => x"2ea63860",
          8125 => x"5902be05",
          8126 => x"22797082",
          8127 => x"055b2378",
          8128 => x"41b43dfe",
          8129 => x"f01153ff",
          8130 => x"840551fe",
          8131 => x"fdbd3f81",
          8132 => x"dccc08df",
          8133 => x"38f7cd39",
          8134 => x"60702254",
          8135 => x"5281d6f8",
          8136 => x"51fef9c0",
          8137 => x"3f80f852",
          8138 => x"7951fefa",
          8139 => x"913f7945",
          8140 => x"79335978",
          8141 => x"ae2ef7ac",
          8142 => x"38789f26",
          8143 => x"87386082",
          8144 => x"0541d539",
          8145 => x"b43dfef0",
          8146 => x"1153ff84",
          8147 => x"0551fefc",
          8148 => x"fa3f81dc",
          8149 => x"cc08802e",
          8150 => x"92386059",
          8151 => x"02be0522",
          8152 => x"79708205",
          8153 => x"5b237841",
          8154 => x"ffae3981",
          8155 => x"d6f051fe",
          8156 => x"f38e3fff",
          8157 => x"a339b43d",
          8158 => x"fef41153",
          8159 => x"ff840551",
          8160 => x"fefcc83f",
          8161 => x"81dccc08",
          8162 => x"802ef6d8",
          8163 => x"38b43dfe",
          8164 => x"f01153ff",
          8165 => x"840551fe",
          8166 => x"fcb13f81",
          8167 => x"dccc0880",
          8168 => x"2ea13860",
          8169 => x"60710c59",
          8170 => x"60840541",
          8171 => x"b43dfef0",
          8172 => x"1153ff84",
          8173 => x"0551fefc",
          8174 => x"923f81dc",
          8175 => x"cc08e438",
          8176 => x"f6a23960",
          8177 => x"70085452",
          8178 => x"81d78451",
          8179 => x"fef8953f",
          8180 => x"80f85279",
          8181 => x"51fef8e6",
          8182 => x"3f794579",
          8183 => x"335978ae",
          8184 => x"2ef68138",
          8185 => x"9f79279c",
          8186 => x"38b43dfe",
          8187 => x"f01153ff",
          8188 => x"840551fe",
          8189 => x"fbd53f81",
          8190 => x"dccc0880",
          8191 => x"2e8d3860",
          8192 => x"60710c59",
          8193 => x"60840541",
          8194 => x"ffb93981",
          8195 => x"d6f051fe",
          8196 => x"f1ee3fff",
          8197 => x"ae39b43d",
          8198 => x"ff801153",
          8199 => x"ff840551",
          8200 => x"fef9b63f",
          8201 => x"81dccc08",
          8202 => x"802ef5b8",
          8203 => x"38635281",
          8204 => x"d79051fe",
          8205 => x"f7ae3f63",
          8206 => x"597804b4",
          8207 => x"3dff8011",
          8208 => x"53ff8405",
          8209 => x"51fef991",
          8210 => x"3f81dccc",
          8211 => x"08802ef5",
          8212 => x"93386352",
          8213 => x"81d7ac51",
          8214 => x"fef7893f",
          8215 => x"6359782d",
          8216 => x"81dccc08",
          8217 => x"802ef4fc",
          8218 => x"3881dccc",
          8219 => x"085281d7",
          8220 => x"c851fef6",
          8221 => x"ef3ff4ec",
          8222 => x"3981d7e4",
          8223 => x"51fef180",
          8224 => x"3ffed5d6",
          8225 => x"3ff4dd39",
          8226 => x"81d88051",
          8227 => x"fef0f13f",
          8228 => x"8059ffa5",
          8229 => x"39feeb9a",
          8230 => x"3ff4c939",
          8231 => x"64703351",
          8232 => x"5978802e",
          8233 => x"f4be387d",
          8234 => x"7d065978",
          8235 => x"802e81d8",
          8236 => x"38b43dff",
          8237 => x"840551fe",
          8238 => x"de993f81",
          8239 => x"dccc085c",
          8240 => x"815b7a82",
          8241 => x"2eb2387a",
          8242 => x"82248938",
          8243 => x"7a812e8c",
          8244 => x"3880cd39",
          8245 => x"7a832eb0",
          8246 => x"3880c539",
          8247 => x"81d89456",
          8248 => x"7b5581d8",
          8249 => x"98548053",
          8250 => x"81d89c52",
          8251 => x"b43dffb0",
          8252 => x"0551fef6",
          8253 => x"853fbb39",
          8254 => x"81d8bc52",
          8255 => x"b43dffb0",
          8256 => x"0551fef5",
          8257 => x"f53fab39",
          8258 => x"7b5581d8",
          8259 => x"98548053",
          8260 => x"81d8ac52",
          8261 => x"b43dffb0",
          8262 => x"0551fef5",
          8263 => x"dd3f9339",
          8264 => x"7b548053",
          8265 => x"81d8b852",
          8266 => x"b43dffb0",
          8267 => x"0551fef5",
          8268 => x"c93f81d8",
          8269 => x"f85881dd",
          8270 => x"80578056",
          8271 => x"64811146",
          8272 => x"81055580",
          8273 => x"54838080",
          8274 => x"53838080",
          8275 => x"52b43dff",
          8276 => x"b00551eb",
          8277 => x"8a3f81dc",
          8278 => x"cc0881dc",
          8279 => x"cc080970",
          8280 => x"30707207",
          8281 => x"8025515b",
          8282 => x"5b5f805a",
          8283 => x"7a832683",
          8284 => x"38815a78",
          8285 => x"7a065978",
          8286 => x"802e8d38",
          8287 => x"811b7081",
          8288 => x"ff065c59",
          8289 => x"7afebb38",
          8290 => x"7d81327d",
          8291 => x"81320759",
          8292 => x"788a387e",
          8293 => x"ff2e0981",
          8294 => x"06f2c938",
          8295 => x"81d8c051",
          8296 => x"fef4c13f",
          8297 => x"f2be39fc",
          8298 => x"3d0d800b",
          8299 => x"81dd8034",
          8300 => x"87c0948c",
          8301 => x"70085455",
          8302 => x"87848052",
          8303 => x"7251fed3",
          8304 => x"b83f81dc",
          8305 => x"cc08902b",
          8306 => x"75085553",
          8307 => x"87848052",
          8308 => x"7351fed3",
          8309 => x"a43f7281",
          8310 => x"dccc0807",
          8311 => x"750c87c0",
          8312 => x"949c7008",
          8313 => x"54558784",
          8314 => x"80527251",
          8315 => x"fed38a3f",
          8316 => x"81dccc08",
          8317 => x"902b7508",
          8318 => x"55538784",
          8319 => x"80527351",
          8320 => x"fed2f63f",
          8321 => x"7281dccc",
          8322 => x"0807750c",
          8323 => x"8c80830b",
          8324 => x"87c09484",
          8325 => x"0c8c8083",
          8326 => x"0b87c094",
          8327 => x"940ca3bc",
          8328 => x"0b81dcdc",
          8329 => x"0ca6bd0b",
          8330 => x"81dce00c",
          8331 => x"fee3b73f",
          8332 => x"feecde3f",
          8333 => x"81d8d051",
          8334 => x"feedc53f",
          8335 => x"81d8dc51",
          8336 => x"feedbd3f",
          8337 => x"81b1cd51",
          8338 => x"feecc13f",
          8339 => x"8151ecbe",
          8340 => x"3ff0c13f",
          8341 => x"80040000",
          8342 => x"00ffffff",
          8343 => x"ff00ffff",
          8344 => x"ffff00ff",
          8345 => x"ffffff00",
          8346 => x"00001863",
          8347 => x"00001869",
          8348 => x"0000186f",
          8349 => x"00001875",
          8350 => x"0000187b",
          8351 => x"000055d4",
          8352 => x"00005558",
          8353 => x"0000555f",
          8354 => x"00005566",
          8355 => x"0000556d",
          8356 => x"00005574",
          8357 => x"0000557b",
          8358 => x"00005582",
          8359 => x"00005589",
          8360 => x"00005590",
          8361 => x"00005597",
          8362 => x"0000559e",
          8363 => x"000055a4",
          8364 => x"000055aa",
          8365 => x"000055b0",
          8366 => x"000055b6",
          8367 => x"000055bc",
          8368 => x"000055c2",
          8369 => x"000055c8",
          8370 => x"000055ce",
          8371 => x"25642f25",
          8372 => x"642f2564",
          8373 => x"2025643a",
          8374 => x"25643a25",
          8375 => x"642e2564",
          8376 => x"25640a00",
          8377 => x"536f4320",
          8378 => x"436f6e66",
          8379 => x"69677572",
          8380 => x"6174696f",
          8381 => x"6e000000",
          8382 => x"20286672",
          8383 => x"6f6d2053",
          8384 => x"6f432063",
          8385 => x"6f6e6669",
          8386 => x"67290000",
          8387 => x"3a0a4465",
          8388 => x"76696365",
          8389 => x"7320696d",
          8390 => x"706c656d",
          8391 => x"656e7465",
          8392 => x"643a0a00",
          8393 => x"20202020",
          8394 => x"57422053",
          8395 => x"4452414d",
          8396 => x"20202825",
          8397 => x"3038583a",
          8398 => x"25303858",
          8399 => x"292e0a00",
          8400 => x"20202020",
          8401 => x"53445241",
          8402 => x"4d202020",
          8403 => x"20202825",
          8404 => x"3038583a",
          8405 => x"25303858",
          8406 => x"292e0a00",
          8407 => x"20202020",
          8408 => x"494e534e",
          8409 => x"20425241",
          8410 => x"4d202825",
          8411 => x"3038583a",
          8412 => x"25303858",
          8413 => x"292e0a00",
          8414 => x"20202020",
          8415 => x"4252414d",
          8416 => x"20202020",
          8417 => x"20202825",
          8418 => x"3038583a",
          8419 => x"25303858",
          8420 => x"292e0a00",
          8421 => x"20202020",
          8422 => x"52414d20",
          8423 => x"20202020",
          8424 => x"20202825",
          8425 => x"3038583a",
          8426 => x"25303858",
          8427 => x"292e0a00",
          8428 => x"20202020",
          8429 => x"53442043",
          8430 => x"41524420",
          8431 => x"20202844",
          8432 => x"65766963",
          8433 => x"6573203d",
          8434 => x"25303264",
          8435 => x"292e0a00",
          8436 => x"20202020",
          8437 => x"54494d45",
          8438 => x"52312020",
          8439 => x"20202854",
          8440 => x"696d6572",
          8441 => x"7320203d",
          8442 => x"25303264",
          8443 => x"292e0a00",
          8444 => x"20202020",
          8445 => x"494e5452",
          8446 => x"20435452",
          8447 => x"4c202843",
          8448 => x"68616e6e",
          8449 => x"656c733d",
          8450 => x"25303264",
          8451 => x"292e0a00",
          8452 => x"20202020",
          8453 => x"57495348",
          8454 => x"424f4e45",
          8455 => x"20425553",
          8456 => x"0a000000",
          8457 => x"20202020",
          8458 => x"57422049",
          8459 => x"32430a00",
          8460 => x"20202020",
          8461 => x"494f4354",
          8462 => x"4c0a0000",
          8463 => x"20202020",
          8464 => x"5053320a",
          8465 => x"00000000",
          8466 => x"20202020",
          8467 => x"5350490a",
          8468 => x"00000000",
          8469 => x"41646472",
          8470 => x"65737365",
          8471 => x"733a0a00",
          8472 => x"20202020",
          8473 => x"43505520",
          8474 => x"52657365",
          8475 => x"74205665",
          8476 => x"63746f72",
          8477 => x"20416464",
          8478 => x"72657373",
          8479 => x"203d2025",
          8480 => x"3038580a",
          8481 => x"00000000",
          8482 => x"20202020",
          8483 => x"43505520",
          8484 => x"4d656d6f",
          8485 => x"72792053",
          8486 => x"74617274",
          8487 => x"20416464",
          8488 => x"72657373",
          8489 => x"203d2025",
          8490 => x"3038580a",
          8491 => x"00000000",
          8492 => x"20202020",
          8493 => x"53746163",
          8494 => x"6b205374",
          8495 => x"61727420",
          8496 => x"41646472",
          8497 => x"65737320",
          8498 => x"20202020",
          8499 => x"203d2025",
          8500 => x"3038580a",
          8501 => x"00000000",
          8502 => x"4d697363",
          8503 => x"3a0a0000",
          8504 => x"20202020",
          8505 => x"5a505520",
          8506 => x"49642020",
          8507 => x"20202020",
          8508 => x"20202020",
          8509 => x"20202020",
          8510 => x"20202020",
          8511 => x"203d2025",
          8512 => x"3034580a",
          8513 => x"00000000",
          8514 => x"20202020",
          8515 => x"53797374",
          8516 => x"656d2043",
          8517 => x"6c6f636b",
          8518 => x"20467265",
          8519 => x"71202020",
          8520 => x"20202020",
          8521 => x"203d2025",
          8522 => x"642e2530",
          8523 => x"34644d48",
          8524 => x"7a0a0000",
          8525 => x"20202020",
          8526 => x"53445241",
          8527 => x"4d20436c",
          8528 => x"6f636b20",
          8529 => x"46726571",
          8530 => x"20202020",
          8531 => x"20202020",
          8532 => x"203d2025",
          8533 => x"642e2530",
          8534 => x"34644d48",
          8535 => x"7a0a0000",
          8536 => x"20202020",
          8537 => x"57697368",
          8538 => x"626f6e65",
          8539 => x"20534452",
          8540 => x"414d2043",
          8541 => x"6c6f636b",
          8542 => x"20467265",
          8543 => x"713d2025",
          8544 => x"642e2530",
          8545 => x"34644d48",
          8546 => x"7a0a0000",
          8547 => x"536d616c",
          8548 => x"6c000000",
          8549 => x"4d656469",
          8550 => x"756d0000",
          8551 => x"466c6578",
          8552 => x"00000000",
          8553 => x"45564f00",
          8554 => x"45564f6d",
          8555 => x"696e0000",
          8556 => x"556e6b6e",
          8557 => x"6f776e00",
          8558 => x"53440000",
          8559 => x"222a2b2c",
          8560 => x"3a3b3c3d",
          8561 => x"3e3f5b5d",
          8562 => x"7c7f0000",
          8563 => x"46415400",
          8564 => x"46415433",
          8565 => x"32000000",
          8566 => x"ebfe904d",
          8567 => x"53444f53",
          8568 => x"352e3000",
          8569 => x"4e4f204e",
          8570 => x"414d4520",
          8571 => x"20202046",
          8572 => x"41543332",
          8573 => x"20202000",
          8574 => x"4e4f204e",
          8575 => x"414d4520",
          8576 => x"20202046",
          8577 => x"41542020",
          8578 => x"20202000",
          8579 => x"000065b8",
          8580 => x"00000000",
          8581 => x"00000000",
          8582 => x"00000000",
          8583 => x"809a4541",
          8584 => x"8e418f80",
          8585 => x"45454549",
          8586 => x"49498e8f",
          8587 => x"9092924f",
          8588 => x"994f5555",
          8589 => x"59999a9b",
          8590 => x"9c9d9e9f",
          8591 => x"41494f55",
          8592 => x"a5a5a6a7",
          8593 => x"a8a9aaab",
          8594 => x"acadaeaf",
          8595 => x"b0b1b2b3",
          8596 => x"b4b5b6b7",
          8597 => x"b8b9babb",
          8598 => x"bcbdbebf",
          8599 => x"c0c1c2c3",
          8600 => x"c4c5c6c7",
          8601 => x"c8c9cacb",
          8602 => x"cccdcecf",
          8603 => x"d0d1d2d3",
          8604 => x"d4d5d6d7",
          8605 => x"d8d9dadb",
          8606 => x"dcdddedf",
          8607 => x"e0e1e2e3",
          8608 => x"e4e5e6e7",
          8609 => x"e8e9eaeb",
          8610 => x"ecedeeef",
          8611 => x"f0f1f2f3",
          8612 => x"f4f5f6f7",
          8613 => x"f8f9fafb",
          8614 => x"fcfdfeff",
          8615 => x"2b2e2c3b",
          8616 => x"3d5b5d2f",
          8617 => x"5c222a3a",
          8618 => x"3c3e3f7c",
          8619 => x"7f000000",
          8620 => x"00010004",
          8621 => x"00100040",
          8622 => x"01000200",
          8623 => x"00000000",
          8624 => x"00010002",
          8625 => x"00040008",
          8626 => x"00100020",
          8627 => x"00000000",
          8628 => x"64696e69",
          8629 => x"74000000",
          8630 => x"64696f63",
          8631 => x"746c0000",
          8632 => x"66696e69",
          8633 => x"74000000",
          8634 => x"666c6f61",
          8635 => x"64000000",
          8636 => x"66657865",
          8637 => x"63000000",
          8638 => x"6d636c65",
          8639 => x"61720000",
          8640 => x"6d636f70",
          8641 => x"79000000",
          8642 => x"6d646966",
          8643 => x"66000000",
          8644 => x"6d64756d",
          8645 => x"70000000",
          8646 => x"6d656200",
          8647 => x"6d656800",
          8648 => x"6d657700",
          8649 => x"68696400",
          8650 => x"68696500",
          8651 => x"68666400",
          8652 => x"68666500",
          8653 => x"63616c6c",
          8654 => x"00000000",
          8655 => x"6a6d7000",
          8656 => x"72657374",
          8657 => x"61727400",
          8658 => x"72657365",
          8659 => x"74000000",
          8660 => x"696e666f",
          8661 => x"00000000",
          8662 => x"74657374",
          8663 => x"00000000",
          8664 => x"74626173",
          8665 => x"69630000",
          8666 => x"4469736b",
          8667 => x"20457272",
          8668 => x"6f720a00",
          8669 => x"496e7465",
          8670 => x"726e616c",
          8671 => x"20657272",
          8672 => x"6f722e0a",
          8673 => x"00000000",
          8674 => x"4469736b",
          8675 => x"206e6f74",
          8676 => x"20726561",
          8677 => x"64792e0a",
          8678 => x"00000000",
          8679 => x"4e6f2066",
          8680 => x"696c6520",
          8681 => x"666f756e",
          8682 => x"642e0a00",
          8683 => x"4e6f2070",
          8684 => x"61746820",
          8685 => x"666f756e",
          8686 => x"642e0a00",
          8687 => x"496e7661",
          8688 => x"6c696420",
          8689 => x"66696c65",
          8690 => x"6e616d65",
          8691 => x"2e0a0000",
          8692 => x"41636365",
          8693 => x"73732064",
          8694 => x"656e6965",
          8695 => x"642e0a00",
          8696 => x"46696c65",
          8697 => x"20616c72",
          8698 => x"65616479",
          8699 => x"20657869",
          8700 => x"7374732e",
          8701 => x"0a000000",
          8702 => x"46696c65",
          8703 => x"2068616e",
          8704 => x"646c6520",
          8705 => x"696e7661",
          8706 => x"6c69642e",
          8707 => x"0a000000",
          8708 => x"53442069",
          8709 => x"73207772",
          8710 => x"69746520",
          8711 => x"70726f74",
          8712 => x"65637465",
          8713 => x"642e0a00",
          8714 => x"44726976",
          8715 => x"65206e75",
          8716 => x"6d626572",
          8717 => x"20697320",
          8718 => x"696e7661",
          8719 => x"6c69642e",
          8720 => x"0a000000",
          8721 => x"4469736b",
          8722 => x"206e6f74",
          8723 => x"20656e61",
          8724 => x"626c6564",
          8725 => x"2e0a0000",
          8726 => x"4e6f2063",
          8727 => x"6f6d7061",
          8728 => x"7469626c",
          8729 => x"65206669",
          8730 => x"6c657379",
          8731 => x"7374656d",
          8732 => x"20666f75",
          8733 => x"6e64206f",
          8734 => x"6e206469",
          8735 => x"736b2e0a",
          8736 => x"00000000",
          8737 => x"466f726d",
          8738 => x"61742061",
          8739 => x"626f7274",
          8740 => x"65642e0a",
          8741 => x"00000000",
          8742 => x"54696d65",
          8743 => x"6f75742c",
          8744 => x"206f7065",
          8745 => x"72617469",
          8746 => x"6f6e2063",
          8747 => x"616e6365",
          8748 => x"6c6c6564",
          8749 => x"2e0a0000",
          8750 => x"46696c65",
          8751 => x"20697320",
          8752 => x"6c6f636b",
          8753 => x"65642e0a",
          8754 => x"00000000",
          8755 => x"496e7375",
          8756 => x"66666963",
          8757 => x"69656e74",
          8758 => x"206d656d",
          8759 => x"6f72792e",
          8760 => x"0a000000",
          8761 => x"546f6f20",
          8762 => x"6d616e79",
          8763 => x"206f7065",
          8764 => x"6e206669",
          8765 => x"6c65732e",
          8766 => x"0a000000",
          8767 => x"50617261",
          8768 => x"6d657465",
          8769 => x"72732069",
          8770 => x"6e636f72",
          8771 => x"72656374",
          8772 => x"2e0a0000",
          8773 => x"53756363",
          8774 => x"6573732e",
          8775 => x"0a000000",
          8776 => x"556e6b6e",
          8777 => x"6f776e20",
          8778 => x"6572726f",
          8779 => x"722e0a00",
          8780 => x"0a256c75",
          8781 => x"20627974",
          8782 => x"65732025",
          8783 => x"73206174",
          8784 => x"20256c75",
          8785 => x"20627974",
          8786 => x"65732f73",
          8787 => x"65632e0a",
          8788 => x"00000000",
          8789 => x"72656164",
          8790 => x"00000000",
          8791 => x"25303858",
          8792 => x"00000000",
          8793 => x"3a202000",
          8794 => x"25303458",
          8795 => x"00000000",
          8796 => x"20202020",
          8797 => x"20202020",
          8798 => x"00000000",
          8799 => x"25303258",
          8800 => x"00000000",
          8801 => x"20200000",
          8802 => x"207c0000",
          8803 => x"7c0d0a00",
          8804 => x"7a4f5300",
          8805 => x"0a2a2a20",
          8806 => x"25732028",
          8807 => x"00000000",
          8808 => x"31302f30",
          8809 => x"342f3230",
          8810 => x"32300000",
          8811 => x"76312e30",
          8812 => x"00000000",
          8813 => x"205a5055",
          8814 => x"2c207265",
          8815 => x"76202530",
          8816 => x"32782920",
          8817 => x"25732025",
          8818 => x"73202a2a",
          8819 => x"0a0a0000",
          8820 => x"5a505520",
          8821 => x"496e7465",
          8822 => x"72727570",
          8823 => x"74204861",
          8824 => x"6e646c65",
          8825 => x"720a0000",
          8826 => x"54696d65",
          8827 => x"7220696e",
          8828 => x"74657272",
          8829 => x"7570740a",
          8830 => x"00000000",
          8831 => x"50533220",
          8832 => x"696e7465",
          8833 => x"72727570",
          8834 => x"740a0000",
          8835 => x"494f4354",
          8836 => x"4c205244",
          8837 => x"20696e74",
          8838 => x"65727275",
          8839 => x"70740a00",
          8840 => x"494f4354",
          8841 => x"4c205752",
          8842 => x"20696e74",
          8843 => x"65727275",
          8844 => x"70740a00",
          8845 => x"55415254",
          8846 => x"30205258",
          8847 => x"20696e74",
          8848 => x"65727275",
          8849 => x"70740a00",
          8850 => x"55415254",
          8851 => x"30205458",
          8852 => x"20696e74",
          8853 => x"65727275",
          8854 => x"70740a00",
          8855 => x"55415254",
          8856 => x"31205258",
          8857 => x"20696e74",
          8858 => x"65727275",
          8859 => x"70740a00",
          8860 => x"55415254",
          8861 => x"31205458",
          8862 => x"20696e74",
          8863 => x"65727275",
          8864 => x"70740a00",
          8865 => x"53657474",
          8866 => x"696e6720",
          8867 => x"75702074",
          8868 => x"696d6572",
          8869 => x"2e2e2e0a",
          8870 => x"00000000",
          8871 => x"456e6162",
          8872 => x"6c696e67",
          8873 => x"2074696d",
          8874 => x"65722e2e",
          8875 => x"2e0a0000",
          8876 => x"6175746f",
          8877 => x"65786563",
          8878 => x"2e626174",
          8879 => x"00000000",
          8880 => x"303a0000",
          8881 => x"4661696c",
          8882 => x"65642074",
          8883 => x"6f20696e",
          8884 => x"69746961",
          8885 => x"6c697365",
          8886 => x"20736420",
          8887 => x"63617264",
          8888 => x"20302c20",
          8889 => x"706c6561",
          8890 => x"73652069",
          8891 => x"6e697420",
          8892 => x"6d616e75",
          8893 => x"616c6c79",
          8894 => x"2e0a0000",
          8895 => x"2a200000",
          8896 => x"436c6561",
          8897 => x"72696e67",
          8898 => x"2e2e2e2e",
          8899 => x"00000000",
          8900 => x"436f7079",
          8901 => x"696e672e",
          8902 => x"2e2e0000",
          8903 => x"436f6d70",
          8904 => x"6172696e",
          8905 => x"672e2e2e",
          8906 => x"00000000",
          8907 => x"2530386c",
          8908 => x"78282530",
          8909 => x"3878292d",
          8910 => x"3e253038",
          8911 => x"6c782825",
          8912 => x"30387829",
          8913 => x"0a000000",
          8914 => x"44756d70",
          8915 => x"204d656d",
          8916 => x"6f72790a",
          8917 => x"00000000",
          8918 => x"0a436f6d",
          8919 => x"706c6574",
          8920 => x"652e0a00",
          8921 => x"25303858",
          8922 => x"20253032",
          8923 => x"582d0000",
          8924 => x"3f3f3f0a",
          8925 => x"00000000",
          8926 => x"25303858",
          8927 => x"20253034",
          8928 => x"582d0000",
          8929 => x"25303858",
          8930 => x"20253038",
          8931 => x"582d0000",
          8932 => x"45786563",
          8933 => x"7574696e",
          8934 => x"6720636f",
          8935 => x"64652040",
          8936 => x"20253038",
          8937 => x"78202e2e",
          8938 => x"2e0a0000",
          8939 => x"43616c6c",
          8940 => x"696e6720",
          8941 => x"636f6465",
          8942 => x"20402025",
          8943 => x"30387820",
          8944 => x"2e2e2e0a",
          8945 => x"00000000",
          8946 => x"43616c6c",
          8947 => x"20726574",
          8948 => x"75726e65",
          8949 => x"6420636f",
          8950 => x"64652028",
          8951 => x"2564292e",
          8952 => x"0a000000",
          8953 => x"52657374",
          8954 => x"61727469",
          8955 => x"6e672061",
          8956 => x"70706c69",
          8957 => x"63617469",
          8958 => x"6f6e2e2e",
          8959 => x"2e0a0000",
          8960 => x"436f6c64",
          8961 => x"20726562",
          8962 => x"6f6f7469",
          8963 => x"6e672e2e",
          8964 => x"2e0a0000",
          8965 => x"5a505500",
          8966 => x"62696e00",
          8967 => x"25643a5c",
          8968 => x"25735c25",
          8969 => x"732e2573",
          8970 => x"00000000",
          8971 => x"25643a5c",
          8972 => x"25735c25",
          8973 => x"73000000",
          8974 => x"25643a5c",
          8975 => x"25730000",
          8976 => x"42616420",
          8977 => x"636f6d6d",
          8978 => x"616e642e",
          8979 => x"0a000000",
          8980 => x"52756e6e",
          8981 => x"696e672e",
          8982 => x"2e2e0a00",
          8983 => x"456e6162",
          8984 => x"6c696e67",
          8985 => x"20696e74",
          8986 => x"65727275",
          8987 => x"7074732e",
          8988 => x"2e2e0a00",
          8989 => x"00000000",
          8990 => x"00000000",
          8991 => x"00007fff",
          8992 => x"00000000",
          8993 => x"00007fff",
          8994 => x"00010000",
          8995 => x"00007fff",
          8996 => x"00010000",
          8997 => x"00810000",
          8998 => x"01000000",
          8999 => x"017fffff",
          9000 => x"00000000",
          9001 => x"00000000",
          9002 => x"00007800",
          9003 => x"00000000",
          9004 => x"05f5e100",
          9005 => x"05f5e100",
          9006 => x"05f5e100",
          9007 => x"00000000",
          9008 => x"01010101",
          9009 => x"01010101",
          9010 => x"01011001",
          9011 => x"01000000",
          9012 => x"00000000",
          9013 => x"01000000",
          9014 => x"00000000",
          9015 => x"000066d0",
          9016 => x"01020100",
          9017 => x"00000000",
          9018 => x"00000000",
          9019 => x"000066d8",
          9020 => x"01040100",
          9021 => x"00000000",
          9022 => x"00000000",
          9023 => x"000066e0",
          9024 => x"01140300",
          9025 => x"00000000",
          9026 => x"00000000",
          9027 => x"000066e8",
          9028 => x"012b0300",
          9029 => x"00000000",
          9030 => x"00000000",
          9031 => x"000066f0",
          9032 => x"01300300",
          9033 => x"00000000",
          9034 => x"00000000",
          9035 => x"000066f8",
          9036 => x"013c0400",
          9037 => x"00000000",
          9038 => x"00000000",
          9039 => x"00006700",
          9040 => x"013d0400",
          9041 => x"00000000",
          9042 => x"00000000",
          9043 => x"00006708",
          9044 => x"013f0400",
          9045 => x"00000000",
          9046 => x"00000000",
          9047 => x"00006710",
          9048 => x"01400400",
          9049 => x"00000000",
          9050 => x"00000000",
          9051 => x"00006718",
          9052 => x"01410400",
          9053 => x"00000000",
          9054 => x"00000000",
          9055 => x"0000671c",
          9056 => x"01420400",
          9057 => x"00000000",
          9058 => x"00000000",
          9059 => x"00006720",
          9060 => x"01430400",
          9061 => x"00000000",
          9062 => x"00000000",
          9063 => x"00006724",
          9064 => x"01500500",
          9065 => x"00000000",
          9066 => x"00000000",
          9067 => x"00006728",
          9068 => x"01510500",
          9069 => x"00000000",
          9070 => x"00000000",
          9071 => x"0000672c",
          9072 => x"01540500",
          9073 => x"00000000",
          9074 => x"00000000",
          9075 => x"00006730",
          9076 => x"01550500",
          9077 => x"00000000",
          9078 => x"00000000",
          9079 => x"00006734",
          9080 => x"01790700",
          9081 => x"00000000",
          9082 => x"00000000",
          9083 => x"0000673c",
          9084 => x"01780700",
          9085 => x"00000000",
          9086 => x"00000000",
          9087 => x"00006740",
          9088 => x"01820800",
          9089 => x"00000000",
          9090 => x"00000000",
          9091 => x"00006748",
          9092 => x"01830800",
          9093 => x"00000000",
          9094 => x"00000000",
          9095 => x"00006750",
          9096 => x"01850800",
          9097 => x"00000000",
          9098 => x"00000000",
          9099 => x"00006758",
          9100 => x"01870800",
          9101 => x"00000000",
          9102 => x"00000000",
          9103 => x"00006760",
          9104 => x"018c0900",
          9105 => x"00000000",
          9106 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

